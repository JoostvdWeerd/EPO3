configuration display_synthesised_cfg of display is
   for synthesised
   end for;
end display_synthesised_cfg;
