configuration colour_behaviour_cfg of colour is
   for behaviour
   end for;
end colour_behaviour_cfg;
