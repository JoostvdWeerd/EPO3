configuration enemy_behaviour_cfg of enemy is
   for behaviour
   end for;
end enemy_behaviour_cfg;
