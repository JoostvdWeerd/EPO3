configuration player_behaviour_cfg of player is
   for behaviour
   end for;
end player_behaviour_cfg;
