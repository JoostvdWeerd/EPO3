configuration display_tb_behaviour_cfg of display_tb is
   for behaviour
      for all: display use configuration work.display_behaviour_cfg;
      end for;
   end for;
end display_tb_behaviour_cfg;
