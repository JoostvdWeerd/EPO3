configuration top_level_synthesised_cfg2 of top_level is
   for synthesised
      for all: counter_two use configuration work.counter_two_behaviour_counter_two_cfg;
      end for;
   end for;
end top_level_synthesised_cfg2;
