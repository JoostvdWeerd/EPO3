
library ieee;
use ieee.std_logic_1164.all;
--library tcb018gbwp7t;
--use tcb018gbwp7t.all;

architecture routed of top_level is

  component BUFFD3BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD3BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL0BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL01BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD0BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD10BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DFQD1BWP7T
    port(CP, D : in std_logic; Q : out std_logic);
  end component;

  component NR2XD0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component MAOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component IND2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component XNR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component DFND1BWP7T
    port(CPN, D : in std_logic; Q, QN : out std_logic);
  end component;

  component AO22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component MOAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AN2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component NR2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INR2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component DFKCNQD1BWP7T
    port(CN, CP, D : in std_logic; Q : out std_logic);
  end component;

  component OAI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component ND3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component AOI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component MUX2ND0BWP7T
    port(I0, I1, S : in std_logic; ZN : out std_logic);
  end component;

  component OR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component CKAN2D8BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component INVD1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component AOI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component AOI211D1BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component OR2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component AOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OA21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component NR4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component AOI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component ND4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component AOI211XD0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component OA211D0BWP7T
    port(A1, A2, B, C : in std_logic; Z : out std_logic);
  end component;

  component MAOI222D1BWP7T
    port(A, B, C : in std_logic; ZN : out std_logic);
  end component;

  component AOI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI33D1BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component OAI211D1BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component INR2XD0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component CKND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component IAO21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OAI32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component AO211D0BWP7T
    port(A1, A2, B, C : in std_logic; Z : out std_logic);
  end component;

  component OAI33D1BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component AN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component INR2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component NR3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component AO21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component IND3D1BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component INVD0BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component OAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component IND4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component OA221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component OAI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component OR4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component CKND1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component CKAN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component AN3D1BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component IOA21D1BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component CKND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D1P5BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INR2D2BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component DFD0BWP7T
    port(CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component INVD5BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component INR3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component CKXOR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component DFKCND1BWP7T
    port(CN, CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  signal FE_PHN16_L1_n_23, FE_PHN15_L1_n_33, FE_PHN14_L1_n_24, FE_PHN13_L1_n_22, FE_PHN12_L1_n_28 : std_logic;
  signal FE_PHN11_L1_n_27, FE_PHN10_L1_n_20, FE_PHN9_L1_n_25, FE_PHN8_L1_n_19, FE_PHN7_L1_n_31 : std_logic;
  signal FE_PHN6_L1_n_30, FE_PHN5_L1_n_29, FE_PHN4_L1_n_21, FE_PHN3_L1_n_34, FE_PHN2_L1_n_32 : std_logic;
  signal FE_PHN1_L1_n_26, FE_OFN0_reset, CTS_6 : std_logic;
  signal count_1_s : std_logic_vector(3 downto 0);
  signal count_2_s : std_logic_vector(3 downto 0);
  signal start_value_s : std_logic_vector(3 downto 0);
  signal L1_range_state_out : std_logic_vector(1 downto 0);
  signal L1_state : std_logic_vector(1 downto 0);
  signal L1_n_0, L1_n_1, L1_n_2, L1_n_3, L1_n_4 : std_logic;
  signal L1_n_5, L1_n_6, L1_n_7, L1_n_8, L1_n_9 : std_logic;
  signal L1_n_10, L1_n_11, L1_n_12, L1_n_13, L1_n_14 : std_logic;
  signal L1_n_15, L1_n_16, L1_n_17, L1_n_18, L1_n_19 : std_logic;
  signal L1_n_20, L1_n_21, L1_n_22, L1_n_23, L1_n_24 : std_logic;
  signal L1_n_25, L1_n_26, L1_n_27, L1_n_28, L1_n_29 : std_logic;
  signal L1_n_30, L1_n_31, L1_n_32, L1_n_33, L1_n_34 : std_logic;
  signal L1_n_35, L1_n_36, L1_n_37, L1_n_38, L1_n_39 : std_logic;
  signal L1_n_40, L1_n_41, L1_n_42, L1_n_43, L1_n_44 : std_logic;
  signal L1_n_45, L1_n_46, L1_n_47, L1_n_48, L1_n_49 : std_logic;
  signal L1_n_50, L1_n_51, L1_n_52, L1_n_53, L1_n_54 : std_logic;
  signal L1_n_55, L1_n_56, L1_n_57, L1_n_58, L1_n_59 : std_logic;
  signal L1_n_60, L1_n_61, L1_n_62, L1_n_63, L1_n_64 : std_logic;
  signal L1_n_65, L1_n_66, L1_n_67, L1_n_68, L1_n_69 : std_logic;
  signal L1_n_70, L1_n_71, L1_n_72, L1_n_73, L1_n_74 : std_logic;
  signal L1_n_75, L1_n_76, L1_n_77, L1_n_78, L1_n_79 : std_logic;
  signal L1_n_80, L1_n_81, L1_n_82, L1_n_83, L1_n_84 : std_logic;
  signal L1_n_85, L1_n_86, L1_n_87, L1_n_88, L1_n_89 : std_logic;
  signal L1_n_90, L1_n_91, L1_n_92, L1_n_93, L1_n_94 : std_logic;
  signal L1_n_95, L1_n_96, L1_n_97, L1_n_98, L1_n_99 : std_logic;
  signal L1_n_100, L1_n_101, L1_n_102, L1_n_103, L1_n_104 : std_logic;
  signal L1_n_105, L1_n_106, L1_n_107, L1_n_108, L1_n_109 : std_logic;
  signal L1_n_110, L1_n_111, L1_n_112, L1_n_113, L1_n_114 : std_logic;
  signal L1_n_115, L1_n_116, L1_n_117, L1_n_118, L1_n_119 : std_logic;
  signal L1_n_120, L1_n_121, L1_n_122, L1_n_123, L1_n_124 : std_logic;
  signal L1_n_125, L1_n_126, L1_n_127, L1_n_128, L1_n_129 : std_logic;
  signal L1_n_130, L1_n_131, L1_n_132, L1_n_133, L1_n_134 : std_logic;
  signal L1_n_135, L1_n_136, L1_n_137, L1_n_138, L1_n_139 : std_logic;
  signal L1_n_140, L1_n_141, L1_n_142, L1_n_143, L1_n_144 : std_logic;
  signal L1_n_145, L1_n_146, L1_n_147, L1_n_148, L1_n_149 : std_logic;
  signal L1_n_150, L1_n_151, L1_n_152, L1_n_153, L1_n_154 : std_logic;
  signal L1_n_155, L1_n_156, L1_n_157, L1_n_158, L1_n_159 : std_logic;
  signal L1_n_160, L1_n_161, L1_n_162, L1_n_163, L1_n_164 : std_logic;
  signal L1_n_165, L1_n_166, L1_n_167, L1_n_168, L1_n_169 : std_logic;
  signal L1_n_170, L1_n_171, L1_n_172, L1_n_173, L1_n_174 : std_logic;
  signal L1_n_175, L1_n_176, L1_n_177, L1_n_178, L1_n_179 : std_logic;
  signal L1_n_180, L1_n_181, L1_n_182, L1_n_183, L1_n_184 : std_logic;
  signal L1_n_185, L1_n_186, L1_n_187, L1_n_188, L1_n_189 : std_logic;
  signal L1_n_190, L1_n_191, L1_n_192, L1_n_193, L1_n_194 : std_logic;
  signal L1_n_195, L1_n_196, L1_n_197, L1_n_198, L1_n_199 : std_logic;
  signal L1_n_200, L1_n_201, L1_n_202, L1_n_203, L1_n_204 : std_logic;
  signal L1_n_205, L1_n_206, L1_n_207, L1_n_208, L1_n_209 : std_logic;
  signal L1_n_210, L1_n_211, L1_n_212, L1_n_213, L1_n_214 : std_logic;
  signal L1_n_215, L1_n_216, L1_n_217, L1_n_218, L1_n_219 : std_logic;
  signal L1_n_220, L1_n_221, L1_n_222, L1_n_223, L1_n_224 : std_logic;
  signal L1_n_225, L1_n_226, L1_n_227, L1_n_228, L1_n_229 : std_logic;
  signal L1_n_230, L1_n_231, L1_n_232, L1_n_233, L1_n_234 : std_logic;
  signal L1_n_235, L1_n_236, L1_n_237, L1_n_238, L1_n_239 : std_logic;
  signal L1_n_240, L1_n_241, L1_n_242, L1_n_243, L1_n_244 : std_logic;
  signal L1_n_245, L1_n_246, L1_n_247, L1_n_248, L1_n_249 : std_logic;
  signal L1_n_250, L1_n_251, L1_n_252, L1_n_253, L1_n_254 : std_logic;
  signal L1_n_255, L1_n_256, L1_n_257, L1_n_258, L1_n_259 : std_logic;
  signal L1_n_260, L1_n_261, L1_n_262, L1_n_263, L1_n_264 : std_logic;
  signal L1_n_265, L1_n_266, L1_n_267, L1_n_268, L1_n_269 : std_logic;
  signal L1_n_270, L1_n_271, L1_n_272, L1_n_273, L1_n_274 : std_logic;
  signal L1_n_275, L1_n_276, L1_n_277, L1_n_278, L1_n_279 : std_logic;
  signal L1_n_280, L1_n_281, L1_n_282, L1_n_283, L1_n_284 : std_logic;
  signal L1_n_285, L1_n_286, L1_n_287, L1_n_288, L1_n_289 : std_logic;
  signal L1_n_290, L1_n_291, L1_n_292, L1_n_293, L1_n_294 : std_logic;
  signal L1_n_295, L1_n_296, L1_n_297, L1_n_298, L1_n_299 : std_logic;
  signal L1_n_300, L1_n_301, L1_n_302, L1_n_303, L1_n_304 : std_logic;
  signal L1_n_305, L1_n_306, L1_n_307, L1_n_308, L1_n_309 : std_logic;
  signal L1_n_310, L1_n_311, L1_n_312, L1_n_313, L1_n_314 : std_logic;
  signal L1_n_315, L1_n_316, L1_n_317, L1_n_318, L1_n_319 : std_logic;
  signal L1_n_320, L1_n_321, L1_n_322, L1_n_323, L1_n_324 : std_logic;
  signal L1_n_325, L1_n_326, L1_n_327, L1_n_328, L1_n_329 : std_logic;
  signal L1_n_330, L1_n_331, L1_n_332, L1_n_333, L1_n_334 : std_logic;
  signal L1_n_335, L1_n_336, L1_n_337, L1_n_338, L1_n_339 : std_logic;
  signal L1_n_340, L1_n_341, L1_n_342, L1_n_343, L1_n_344 : std_logic;
  signal L1_n_345, L1_n_346, L1_n_347, L1_n_348, L1_n_349 : std_logic;
  signal L1_n_350, L1_n_351, L1_n_352, L1_n_353, L1_n_354 : std_logic;
  signal L1_n_355, L1_n_356, L1_n_357, L1_n_358, L1_n_359 : std_logic;
  signal L1_n_360, L1_n_361, L1_n_362, L1_n_363, L1_n_364 : std_logic;
  signal L1_n_365, L1_n_366, L1_n_367, L1_n_368, L1_n_369 : std_logic;
  signal L1_n_370, L1_n_371, L1_n_372, L1_n_373, L1_n_374 : std_logic;
  signal L1_n_375, L1_n_376, L1_n_377, L1_n_378, L1_n_379 : std_logic;
  signal L1_n_380, L1_n_381, L1_n_382, L1_n_383, L1_n_384 : std_logic;
  signal L1_n_385, L1_n_386, L1_n_387, L1_n_388, L1_n_389 : std_logic;
  signal L1_n_390, L1_n_391, L1_n_392, L1_n_393, L1_n_394 : std_logic;
  signal L1_n_395, L1_n_396, L1_n_397, L1_n_398, L1_n_399 : std_logic;
  signal L1_n_400, L1_n_401, L1_n_402, L1_n_403, L1_n_404 : std_logic;
  signal L1_n_405, L1_n_406, L1_n_407, L1_n_408, L1_n_409 : std_logic;
  signal L1_n_410, L1_n_411, L1_n_412, L1_n_413, L1_n_414 : std_logic;
  signal L1_n_415, L1_n_416, L1_n_417, L1_n_418, L1_n_419 : std_logic;
  signal L1_n_420, L1_n_421, L1_n_422, L1_n_423, L1_n_424 : std_logic;
  signal L1_n_425, L1_n_426, L1_n_427, L1_n_428, L1_n_429 : std_logic;
  signal L1_n_430, L1_n_431, L1_n_432, L1_n_433, L1_n_434 : std_logic;
  signal L1_n_435, L1_n_436, L1_n_437, L1_n_438, L1_n_439 : std_logic;
  signal L1_n_440, L1_n_441, L1_n_442, L1_n_443, L1_n_444 : std_logic;
  signal L1_n_445, L1_n_446, L1_n_447, L1_n_448, L1_n_449 : std_logic;
  signal L1_n_450, L1_n_451, L1_n_452, L1_n_453, L1_n_454 : std_logic;
  signal L1_n_455, L1_n_456, L1_n_457, L1_n_458, L1_n_459 : std_logic;
  signal L1_n_460, L1_n_461, L1_n_462, L1_n_463, L1_n_464 : std_logic;
  signal L1_n_465, L1_n_466, L1_n_467, L1_n_468, L1_n_469 : std_logic;
  signal L1_n_470, L1_n_471, L1_n_472, L1_n_473, L1_n_474 : std_logic;
  signal L1_n_475, L1_n_476, L1_n_477, L1_n_478, L1_n_479 : std_logic;
  signal L1_n_480, L1_n_481, L1_n_482, L1_n_483, L1_n_484 : std_logic;
  signal L1_n_485, L1_n_486, L1_n_487, L1_n_488, L1_n_489 : std_logic;
  signal L1_n_490, L1_n_491, L1_n_492, L1_n_493, L1_n_494 : std_logic;
  signal L1_n_495, L1_n_496, L1_n_497, L1_n_498, L1_n_499 : std_logic;
  signal L1_n_500, L1_n_501, L1_n_502, L1_n_503, L1_n_504 : std_logic;
  signal L1_n_505, L1_n_506, L1_n_508, L1_n_509, L1_n_510 : std_logic;
  signal L1_n_511, L1_n_512, L1_n_513, L1_n_514, L1_n_515 : std_logic;
  signal L1_n_516, L1_n_517, L1_n_518, L1_n_519, L1_n_520 : std_logic;
  signal L1_n_521, L1_n_522, L1_n_523, L1_n_524, L1_n_525 : std_logic;
  signal L1_n_526, L1_n_527, L1_n_528, L1_n_529, L1_n_530 : std_logic;
  signal L1_n_531, L1_n_532, L1_n_533, L1_n_534, L1_n_535 : std_logic;
  signal L1_n_536, L1_n_537, L1_n_538, L1_n_539, L1_n_540 : std_logic;
  signal L1_n_541, L1_n_542, L1_n_543, L1_n_544, L1_n_545 : std_logic;
  signal L1_n_546, L1_n_547, L1_n_548, L1_n_549, L1_n_550 : std_logic;
  signal L1_n_551, L1_n_552, L1_n_553, L1_n_554, L1_n_555 : std_logic;
  signal L1_n_556, L1_n_557, L1_n_558, L1_n_559, L1_n_560 : std_logic;
  signal L1_n_561, L1_n_562, L1_n_563, L1_n_564, L1_n_565 : std_logic;
  signal L1_n_566, L1_n_567, L1_n_568, L1_n_569, L1_n_570 : std_logic;
  signal L1_n_571, L1_n_573, L1_n_575, L1_n_576, L1_n_577 : std_logic;
  signal L1_n_578, L1_n_579, L1_n_580, L1_n_581, L1_n_582 : std_logic;
  signal L1_n_583, L1_n_584, L1_n_585, L1_n_586, L1_n_587 : std_logic;
  signal L1_n_588, L1_n_589, L1_n_591, L1_n_592, L1_n_594 : std_logic;
  signal L1_n_595, L1_n_596, L1_n_597, L1_n_598, L1_n_599 : std_logic;
  signal L1_n_600, L1_n_601, L1_n_602, L1_n_603, L1_n_604 : std_logic;
  signal L1_n_606, L1_n_608, L1_n_609, L1_n_610, L1_n_611 : std_logic;
  signal L1_n_612, L1_n_613, L1_n_614, L1_n_615, L1_n_616 : std_logic;
  signal L1_n_617, L1_n_618, L1_n_619, L1_n_620, L1_n_621 : std_logic;
  signal L1_n_622, L1_n_623, L1_n_625, L1_n_626, L1_n_627 : std_logic;
  signal L1_n_628, L1_n_629, L1_n_630, L1_n_631, L1_n_632 : std_logic;
  signal L1_n_633, L1_n_634, L1_n_635, L1_n_636, L1_n_637 : std_logic;
  signal L1_n_638, L1_n_639, L1_n_640, L1_n_641, L1_n_642 : std_logic;
  signal L1_n_643, L1_n_644, L1_n_645, L1_n_646, L1_n_647 : std_logic;
  signal L1_n_648, L1_n_649, L1_n_650, L1_n_651, L1_n_652 : std_logic;
  signal L1_n_653, L1_n_654, L1_n_655, L1_n_656, L1_n_657 : std_logic;
  signal L1_n_658, L1_n_659, L1_n_660, L1_n_661, L1_n_662 : std_logic;
  signal L1_n_663, L1_n_664, L1_n_665, L1_n_666, L1_n_667 : std_logic;
  signal L1_n_668, L1_n_669, L1_n_670, L1_n_671, L1_n_672 : std_logic;
  signal L1_n_673, L1_n_674, L1_n_675, L1_n_676, L1_n_677 : std_logic;
  signal L1_n_678, L1_n_679, L1_n_680, L1_n_681, L1_n_682 : std_logic;
  signal L1_n_683, L1_n_684, L1_n_685, L1_n_686, L1_n_688 : std_logic;
  signal L1_n_689, L1_n_691, L1_n_692, L1_n_693, L1_n_694 : std_logic;
  signal L1_n_695, L1_n_696, L1_n_697, L1_n_698, L1_n_699 : std_logic;
  signal L1_n_700, L1_n_701, L1_n_702, L1_n_719, L1_n_723 : std_logic;
  signal L1_n_724, L1_n_725, L1_n_726, L2_n_0, L2_n_1 : std_logic;
  signal L2_n_2, L2_n_3, L2_n_4, L2_n_5, L2_n_6 : std_logic;
  signal L2_n_7, L2_n_8, L2_n_9, L2_n_10, L3_n_0 : std_logic;
  signal L3_n_1, L3_n_2, L3_n_3, L3_n_4, L3_n_5 : std_logic;
  signal L3_n_6, L3_n_7, L3_n_8, L3_n_9, L3_n_10 : std_logic;
  signal L3_n_11, UNCONNECTED, UNCONNECTED0, UNCONNECTED1, enable_s : std_logic;
  signal reset_2_s : std_logic;

begin

  FE_PHC16_L1_n_23 : BUFFD3BWP7T port map(I => L1_n_23, Z => FE_PHN16_L1_n_23);
  FE_PHC15_L1_n_33 : CKBD3BWP7T port map(I => FE_PHN15_L1_n_33, Z => L1_n_33);
  FE_PHC14_L1_n_24 : CKBD3BWP7T port map(I => L1_n_24, Z => FE_PHN14_L1_n_24);
  FE_PHC13_L1_n_22 : DEL0BWP7T port map(I => L1_n_22, Z => FE_PHN13_L1_n_22);
  FE_PHC12_L1_n_28 : DEL01BWP7T port map(I => L1_n_28, Z => FE_PHN12_L1_n_28);
  FE_PHC11_L1_n_27 : DEL01BWP7T port map(I => L1_n_27, Z => FE_PHN11_L1_n_27);
  FE_PHC10_L1_n_20 : DEL01BWP7T port map(I => L1_n_20, Z => FE_PHN10_L1_n_20);
  FE_PHC9_L1_n_25 : DEL01BWP7T port map(I => L1_n_25, Z => FE_PHN9_L1_n_25);
  FE_PHC8_L1_n_19 : DEL01BWP7T port map(I => L1_n_19, Z => FE_PHN8_L1_n_19);
  FE_PHC7_L1_n_31 : DEL01BWP7T port map(I => L1_n_31, Z => FE_PHN7_L1_n_31);
  FE_PHC6_L1_n_30 : DEL01BWP7T port map(I => L1_n_30, Z => FE_PHN6_L1_n_30);
  FE_PHC5_L1_n_29 : CKBD0BWP7T port map(I => L1_n_29, Z => FE_PHN5_L1_n_29);
  FE_PHC4_L1_n_21 : DEL01BWP7T port map(I => L1_n_21, Z => FE_PHN4_L1_n_21);
  FE_PHC3_L1_n_34 : CKBD0BWP7T port map(I => L1_n_34, Z => FE_PHN3_L1_n_34);
  FE_PHC2_L1_n_32 : CKBD0BWP7T port map(I => L1_n_32, Z => FE_PHN2_L1_n_32);
  FE_PHC1_L1_n_26 : CKBD0BWP7T port map(I => L1_n_26, Z => FE_PHN1_L1_n_26);
  FE_OFC0_reset : DEL01BWP7T port map(I => reset, Z => FE_OFN0_reset);
  CTS_ccl_a_BUF_clk_G0_L1_1 : CKBD10BWP7T port map(I => clk, Z => CTS_6);
  L2_count_inside_reg_3 : DFQD1BWP7T port map(CP => CTS_6, D => L2_n_10, Q => count_1_s(3));
  L2_g70 : NR2XD0BWP7T port map(A1 => L2_n_9, A2 => FE_OFN0_reset, ZN => L2_n_10);
  L2_count_inside_reg_2 : DFQD1BWP7T port map(CP => CTS_6, D => L2_n_8, Q => count_1_s(2));
  L2_g72 : MAOI22D0BWP7T port map(A1 => L2_n_5, A2 => count_1_s(3), B1 => L2_n_5, B2 => count_1_s(3), ZN => L2_n_9);
  L2_g73 : NR2XD0BWP7T port map(A1 => L2_n_7, A2 => FE_OFN0_reset, ZN => L2_n_8);
  L2_count_inside_reg_1 : DFQD1BWP7T port map(CP => CTS_6, D => L2_n_6, Q => count_1_s(1));
  L2_g75 : MAOI22D0BWP7T port map(A1 => L2_n_3, A2 => count_1_s(2), B1 => L2_n_3, B2 => count_1_s(2), ZN => L2_n_7);
  L2_g76 : NR2XD0BWP7T port map(A1 => L2_n_4, A2 => FE_OFN0_reset, ZN => L2_n_6);
  L2_g77 : IND2D1BWP7T port map(A1 => L2_n_3, B1 => count_1_s(2), ZN => L2_n_5);
  L2_count_inside_reg_0 : DFQD1BWP7T port map(CP => CTS_6, D => L2_n_2, Q => count_1_s(0));
  L2_g79 : MAOI22D0BWP7T port map(A1 => L2_n_0, A2 => count_1_s(1), B1 => L2_n_0, B2 => count_1_s(1), ZN => L2_n_4);
  L2_g80 : IND2D1BWP7T port map(A1 => L2_n_0, B1 => count_1_s(1), ZN => L2_n_3);
  L2_g81 : NR2XD0BWP7T port map(A1 => L2_n_1, A2 => FE_OFN0_reset, ZN => L2_n_2);
  L2_g82 : XNR2D1BWP7T port map(A1 => enable_s, A2 => count_1_s(0), ZN => L2_n_1);
  L2_g83 : ND2D1BWP7T port map(A1 => enable_s, A2 => count_1_s(0), ZN => L2_n_0);
  L3_count_inside_reg_3 : DFND1BWP7T port map(CPN => CTS_6, D => L3_n_11, Q => count_2_s(3), QN => UNCONNECTED);
  L3_g182 : AO22D0BWP7T port map(A1 => L3_n_9, A2 => L3_n_3, B1 => L3_n_1, B2 => start_value_s(3), Z => L3_n_11);
  L3_count_inside_reg_2 : DFND1BWP7T port map(CPN => CTS_6, D => L3_n_10, Q => count_2_s(2), QN => UNCONNECTED0);
  L3_g184 : AO22D0BWP7T port map(A1 => L3_n_8, A2 => L3_n_3, B1 => L3_n_1, B2 => start_value_s(2), Z => L3_n_10);
  L3_g185 : MOAI22D0BWP7T port map(A1 => L3_n_7, A2 => count_2_s(3), B1 => L3_n_7, B2 => count_2_s(3), ZN => L3_n_9);
  L3_count_inside_reg_1 : DFND1BWP7T port map(CPN => CTS_6, D => L3_n_6, Q => count_2_s(1), QN => UNCONNECTED1);
  L3_g187 : MOAI22D0BWP7T port map(A1 => L3_n_2, A2 => count_2_s(2), B1 => L3_n_2, B2 => count_2_s(2), ZN => L3_n_8);
  L3_count_inside_reg_0 : DFND1BWP7T port map(CPN => CTS_6, D => L3_n_5, Q => count_2_s(0), QN => L3_n_0);
  L3_g189 : AN2D0BWP7T port map(A1 => L3_n_4, A2 => L3_n_3, Z => L3_n_6);
  L3_g190 : IND2D1BWP7T port map(A1 => L3_n_2, B1 => count_2_s(2), ZN => L3_n_7);
  L3_g191 : AO22D0BWP7T port map(A1 => L3_n_0, A2 => L3_n_3, B1 => L3_n_1, B2 => start_value_s(0), Z => L3_n_5);
  L3_g192 : MOAI22D0BWP7T port map(A1 => L3_n_0, A2 => count_2_s(1), B1 => L3_n_0, B2 => count_2_s(1), ZN => L3_n_4);
  L3_g193 : NR2D0BWP7T port map(A1 => reset_2_s, A2 => FE_OFN0_reset, ZN => L3_n_3);
  L3_g194 : ND2D1BWP7T port map(A1 => count_2_s(0), A2 => count_2_s(1), ZN => L3_n_2);
  L3_g195 : INR2D0BWP7T port map(A1 => reset_2_s, B1 => FE_OFN0_reset, ZN => L3_n_1);
  L1_range_state_out_reg_1 : DFKCNQD1BWP7T port map(CN => L1_n_35, CP => CTS_6, D => L1_n_700, Q => L1_range_state_out(1));
  L1_g3348 : OAI221D0BWP7T port map(A1 => L1_n_699, A2 => count_1_s(3), B1 => count_2_s(3), B2 => L1_n_697, C => L1_n_695, ZN => L1_n_701);
  L1_g3349 : ND3D0BWP7T port map(A1 => L1_n_698, A2 => L1_n_696, A3 => L1_n_695, ZN => L1_n_700);
  L1_g3350 : AOI21D0BWP7T port map(A1 => L1_n_696, A2 => count_2_s(3), B => L1_n_691, ZN => L1_n_699);
  L1_g3351 : MOAI22D0BWP7T port map(A1 => L1_n_695, A2 => L1_n_689, B1 => L1_n_689, B2 => count_1_s(2), ZN => start_value_s(2));
  L1_g3352 : MUX2ND0BWP7T port map(I0 => L1_n_693, I1 => L1_n_694, S => count_2_s(3), ZN => L1_n_698);
  L1_g3353 : IND2D1BWP7T port map(A1 => start_value_s(3), B1 => L1_n_694, ZN => start_value_s(0));
  L1_g3354 : IND2D1BWP7T port map(A1 => L1_n_693, B1 => count_2_s(2), ZN => L1_n_697);
  L1_g3355 : IND2D1BWP7T port map(A1 => count_2_s(2), B1 => L1_n_692, ZN => L1_n_696);
  L1_g3356 : OR2D1BWP7T port map(A1 => L1_n_691, A2 => count_1_s(2), Z => L1_n_695);
  L1_g3357 : OR2D1BWP7T port map(A1 => L1_n_691, A2 => count_1_s(3), Z => L1_n_694);
  L1_g3358 : ND2D1BWP7T port map(A1 => L1_n_692, A2 => count_1_s(3), ZN => L1_n_693);
  L1_g3359 : CKAN2D8BWP7T port map(A1 => L1_n_688, A2 => L1_n_18, Z => done);
  L1_g3360 : IND2D1BWP7T port map(A1 => enable_s, B1 => L1_state(0), ZN => reset_2_s);
  L1_g3361 : NR2XD0BWP7T port map(A1 => count_1_s(3), A2 => count_1_s(2), ZN => start_value_s(3));
  L1_g3362 : IND2D1BWP7T port map(A1 => count_1_s(0), B1 => L1_n_689, ZN => L1_n_702);
  L1_g3363 : NR2XD0BWP7T port map(A1 => count_2_s(0), A2 => count_2_s(1), ZN => L1_n_692);
  L1_g3364 : OR2D1BWP7T port map(A1 => count_1_s(0), A2 => count_1_s(1), Z => L1_n_691);
  L1_g3366 : INVD1BWP7T port map(I => count_1_s(3), ZN => L1_n_689);
  L1_state_reg_0 : DFND1BWP7T port map(CPN => CTS_6, D => L1_n_686, Q => L1_state(0), QN => L1_n_18);
  L1_state_reg_1 : DFND1BWP7T port map(CPN => CTS_6, D => L1_n_685, Q => enable_s, QN => L1_n_688);
  L1_g28933 : AOI31D0BWP7T port map(A1 => L1_n_684, A2 => L1_n_145, A3 => L1_n_74, B => FE_OFN0_reset, ZN => L1_n_686);
  L1_g28935 : AOI211D1BWP7T port map(A1 => L1_n_682, A2 => L1_n_98, B => reset_2_s, C => FE_OFN0_reset, ZN => L1_n_685);
  L1_g28936 : OR2D0BWP7T port map(A1 => L1_n_683, A2 => enable_s, Z => L1_n_684);
  L1_g28937 : AOI22D0BWP7T port map(A1 => L1_n_681, A2 => L1_state(0), B1 => L1_n_18, B2 => main_enable, ZN => L1_n_683);
  L1_g28938 : OA21D0BWP7T port map(A1 => L1_n_45, A2 => start_value_s(0), B => L1_n_681, Z => L1_n_682);
  L1_g28939 : NR4D0BWP7T port map(A1 => L1_n_680, A2 => L1_n_655, A3 => L1_n_633, A4 => L1_n_609, ZN => L1_n_681);
  L1_g28940 : AOI221D0BWP7T port map(A1 => L1_n_719, A2 => L1_n_526, B1 => L1_n_726, B2 => L1_n_525, C => L1_n_679, ZN => L1_n_680);
  L1_g28941 : ND4D0BWP7T port map(A1 => L1_n_678, A2 => L1_n_672, A3 => L1_n_676, A4 => L1_n_315, ZN => L1_n_679);
  L1_g28942 : AOI211XD0BWP7T port map(A1 => L1_n_662, A2 => L1_n_524, B => L1_n_675, C => L1_n_677, ZN => L1_n_678);
  L1_g28943 : OA211D0BWP7T port map(A1 => L1_n_524, A2 => L1_n_662, B => L1_n_674, C => L1_n_673, Z => L1_n_677);
  L1_g28944 : OAI221D0BWP7T port map(A1 => L1_n_726, A2 => L1_n_525, B1 => L1_n_496, B2 => L1_n_659, C => L1_n_669, ZN => L1_n_676);
  L1_g28945 : MAOI222D1BWP7T port map(A => L1_n_670, B => L1_n_640, C => L1_n_526, ZN => L1_n_675);
  L1_g28946 : AOI222D0BWP7T port map(A1 => L1_n_671, A2 => L1_n_527, B1 => L1_n_668, B2 => L1_n_644, C1 => L1_n_647, C2 => L1_n_522, ZN => L1_n_674);
  L1_g28947 : AOI33D1BWP7T port map(A1 => L1_n_663, A2 => L1_n_598, A3 => L1_n_520, B1 => L1_n_660, B2 => L1_n_626, B3 => L1_n_496, ZN => L1_n_673);
  L1_g28948 : OAI211D1BWP7T port map(A1 => L1_n_526, A2 => L1_n_719, B => L1_n_667, C => L1_n_658, ZN => L1_n_672);
  L1_g28949 : INR2XD0BWP7T port map(A1 => L1_n_668, B1 => L1_n_603, ZN => L1_n_671);
  L1_g28950 : CKND2D1BWP7T port map(A1 => L1_n_665, A2 => L1_n_666, ZN => L1_n_670);
  L1_g28951 : AOI21D0BWP7T port map(A1 => L1_n_657, A2 => L1_n_639, B => L1_n_664, ZN => L1_n_669);
  L1_g28952 : AOI221D0BWP7T port map(A1 => L1_n_652, A2 => L1_n_646, B1 => L1_n_642, B2 => L1_n_493, C => L1_n_650, ZN => L1_n_667);
  L1_g28953 : OA21D0BWP7T port map(A1 => L1_n_598, A2 => L1_n_520, B => L1_n_663, Z => L1_n_668);
  L1_g28954 : AOI31D0BWP7T port map(A1 => L1_n_648, A2 => L1_n_608, A3 => L1_n_503, B => L1_n_661, ZN => L1_n_666);
  L1_g28955 : AOI33D1BWP7T port map(A1 => L1_n_653, A2 => L1_n_617, A3 => L1_n_502, B1 => L1_n_643, B2 => L1_n_630, B3 => L1_n_497, ZN => L1_n_665);
  L1_g28956 : MOAI22D0BWP7T port map(A1 => L1_n_645, A2 => L1_n_522, B1 => L1_n_657, B2 => L1_n_651, ZN => L1_n_664);
  L1_g28957 : OA21D0BWP7T port map(A1 => L1_n_626, A2 => L1_n_496, B => L1_n_660, Z => L1_n_663);
  L1_g28958 : OAI21D0BWP7T port map(A1 => L1_n_629, A2 => L1_n_493, B => L1_n_656, ZN => L1_n_661);
  L1_g28959 : MAOI22D0BWP7T port map(A1 => L1_n_641, A2 => L1_n_517, B1 => L1_n_641, B2 => L1_n_517, ZN => L1_n_662);
  L1_g28960 : ND2D1BWP7T port map(A1 => L1_n_654, A2 => L1_n_625, ZN => L1_n_659);
  L1_g28961 : ND2D1BWP7T port map(A1 => L1_n_649, A2 => L1_n_646, ZN => L1_n_658);
  L1_g28962 : OR2D1BWP7T port map(A1 => L1_n_647, A2 => L1_n_522, Z => L1_n_660);
  L1_g28963 : OAI211D1BWP7T port map(A1 => L1_n_502, A2 => L1_n_617, B => L1_n_653, C => L1_n_638, ZN => L1_n_656);
  L1_g28964 : AOI211XD0BWP7T port map(A1 => L1_n_637, A2 => L1_n_632, B => L1_n_627, C => L1_n_719, ZN => L1_n_655);
  L1_g28965 : OA21D0BWP7T port map(A1 => L1_n_625, A2 => L1_n_495, B => L1_n_654, Z => L1_n_657);
  L1_g28966 : AOI211XD0BWP7T port map(A1 => L1_n_612, A2 => L1_n_502, B => L1_n_635, C => L1_n_634, ZN => L1_n_652);
  L1_g28967 : ND2D1BWP7T port map(A1 => L1_n_645, A2 => L1_n_522, ZN => L1_n_654);
  L1_g28968 : OA21D0BWP7T port map(A1 => L1_n_608, A2 => L1_n_503, B => L1_n_648, Z => L1_n_653);
  L1_g28969 : AOI211XD0BWP7T port map(A1 => L1_n_616, A2 => L1_n_527, B => L1_n_636, C => L1_n_620, ZN => L1_n_651);
  L1_g28970 : IAO21D0BWP7T port map(A1 => L1_n_642, A2 => L1_n_493, B => L1_n_627, ZN => L1_n_650);
  L1_g28971 : OAI32D1BWP7T port map(A1 => L1_n_502, A2 => L1_n_612, A3 => L1_n_634, B1 => L1_n_503, B2 => L1_n_628, ZN => L1_n_649);
  L1_g28972 : OA21D0BWP7T port map(A1 => L1_n_630, A2 => L1_n_497, B => L1_n_643, Z => L1_n_648);
  L1_g28973 : AOI21D0BWP7T port map(A1 => L1_n_618, A2 => L1_n_513, B => L1_n_641, ZN => L1_n_647);
  L1_g28974 : AOI211XD0BWP7T port map(A1 => L1_n_582, A2 => L1_n_521, B => L1_n_631, C => L1_n_610, ZN => L1_n_644);
  L1_g28975 : AOI22D0BWP7T port map(A1 => L1_n_627, A2 => L1_n_492, B1 => L1_n_632, B2 => L1_n_497, ZN => L1_n_646);
  L1_g28976 : MAOI22D0BWP7T port map(A1 => L1_n_619, A2 => L1_n_513, B1 => L1_n_619, B2 => L1_n_513, ZN => L1_n_645);
  L1_g28977 : ND2D1BWP7T port map(A1 => L1_n_629, A2 => L1_n_493, ZN => L1_n_643);
  L1_g28978 : ND2D1BWP7T port map(A1 => L1_n_621, A2 => L1_n_532, ZN => L1_n_640);
  L1_g28979 : NR2XD0BWP7T port map(A1 => L1_n_632, A2 => L1_n_497, ZN => L1_n_642);
  L1_g28980 : NR2D1BWP7T port map(A1 => L1_n_618, A2 => L1_n_513, ZN => L1_n_641);
  L1_g28981 : OAI32D1BWP7T port map(A1 => L1_n_527, A2 => L1_n_616, A3 => L1_n_620, B1 => L1_n_520, B2 => L1_n_595, ZN => L1_n_639);
  L1_g28982 : MAOI222D1BWP7T port map(A => L1_n_615, B => L1_n_579, C => L1_n_505, ZN => L1_n_638);
  L1_g28983 : AO211D0BWP7T port map(A1 => L1_n_604, A2 => L1_n_596, B => L1_n_628, C => L1_n_612, Z => L1_n_637);
  L1_g28984 : MAOI222D1BWP7T port map(A => L1_n_622, B => L1_n_723, C => L1_n_521, ZN => L1_n_636);
  L1_g28985 : MAOI222D1BWP7T port map(A => L1_n_614, B => L1_n_597, C => L1_n_505, ZN => L1_n_635);
  L1_g28986 : OAI33D1BWP7T port map(A1 => L1_n_514, A2 => L1_n_512, A3 => L1_n_606, B1 => L1_n_489, B2 => L1_n_542, B3 => L1_n_586, ZN => L1_n_633);
  L1_g28987 : AN2D1BWP7T port map(A1 => L1_n_628, A2 => L1_n_503, Z => L1_n_634);
  L1_g28988 : OA21D0BWP7T port map(A1 => L1_n_582, A2 => L1_n_521, B => L1_n_623, Z => L1_n_631);
  L1_g28989 : MAOI22D0BWP7T port map(A1 => L1_n_602, A2 => L1_n_514, B1 => L1_n_602, B2 => L1_n_514, ZN => L1_n_632);
  L1_g28990 : AOI211XD0BWP7T port map(A1 => L1_n_581, A2 => L1_n_514, B => L1_n_613, C => L1_n_534, ZN => L1_n_630);
  L1_g28991 : OAI21D0BWP7T port map(A1 => L1_n_613, A2 => L1_n_511, B => L1_n_621, ZN => L1_n_629);
  L1_g28992 : AOI211D1BWP7T port map(A1 => L1_n_587, A2 => L1_n_484, B => L1_n_600, C => L1_n_71, ZN => L1_n_628);
  L1_g28993 : AOI211D1BWP7T port map(A1 => L1_n_601, A2 => L1_n_512, B => L1_n_611, C => L1_n_71, ZN => L1_n_627);
  L1_g28994 : MAOI222D1BWP7T port map(A => L1_n_599, B => L1_n_576, C => L1_n_523, ZN => L1_n_623);
  L1_g28995 : MAOI222D1BWP7T port map(A => L1_n_592, B => L1_n_584, C => L1_n_523, ZN => L1_n_622);
  L1_g28996 : OA21D0BWP7T port map(A1 => L1_n_589, A2 => L1_n_509, B => L1_n_618, Z => L1_n_626);
  L1_g28997 : MOAI22D0BWP7T port map(A1 => L1_n_588, A2 => L1_n_510, B1 => L1_n_588, B2 => L1_n_510, ZN => L1_n_625);
  L1_g28999 : ND2D1BWP7T port map(A1 => L1_n_613, A2 => L1_n_511, ZN => L1_n_621);
  L1_g29000 : AN2D1BWP7T port map(A1 => L1_n_595, A2 => L1_n_520, Z => L1_n_620);
  L1_g29001 : OR2D1BWP7T port map(A1 => L1_n_588, A2 => L1_n_509, Z => L1_n_619);
  L1_g29002 : ND2D1BWP7T port map(A1 => L1_n_589, A2 => L1_n_509, ZN => L1_n_618);
  L1_g29003 : MOAI22D0BWP7T port map(A1 => L1_n_564, A2 => L1_n_531, B1 => L1_n_564, B2 => L1_n_531, ZN => L1_n_617);
  L1_g29004 : MAOI22D0BWP7T port map(A1 => L1_n_570, A2 => L1_n_518, B1 => L1_n_570, B2 => L1_n_518, ZN => L1_n_616);
  L1_g29005 : MAOI22D0BWP7T port map(A1 => L1_n_567, A2 => L1_n_498, B1 => L1_n_594, B2 => L1_n_585, ZN => L1_n_615);
  L1_g29006 : MAOI222D1BWP7T port map(A => L1_n_573, B => L1_n_591, C => L1_n_498, ZN => L1_n_614);
  L1_g29007 : NR2XD0BWP7T port map(A1 => L1_n_601, A2 => L1_n_512, ZN => L1_n_611);
  L1_g29008 : INR2D1BWP7T port map(A1 => L1_n_603, B1 => L1_n_527, ZN => L1_n_610);
  L1_g29009 : AOI21D0BWP7T port map(A1 => L1_n_578, A2 => L1_n_540, B => L1_n_516, ZN => L1_n_609);
  L1_g29010 : NR3D0BWP7T port map(A1 => L1_n_581, A2 => L1_n_485, A3 => L1_n_514, ZN => L1_n_613);
  L1_g29011 : AOI211D1BWP7T port map(A1 => L1_n_566, A2 => L1_n_531, B => L1_n_583, C => L1_n_71, ZN => L1_n_612);
  L1_g29012 : AO21D0BWP7T port map(A1 => L1_n_575, A2 => L1_n_485, B => L1_n_532, Z => L1_n_606);
  L1_g29014 : IND3D1BWP7T port map(A1 => L1_n_591, B1 => L1_n_499, B2 => L1_n_555, ZN => L1_n_604);
  L1_g29015 : MOAI22D0BWP7T port map(A1 => L1_n_581, A2 => L1_n_484, B1 => L1_n_581, B2 => L1_n_484, ZN => L1_n_608);
  L1_g29017 : NR2XD0BWP7T port map(A1 => L1_n_587, A2 => L1_n_484, ZN => L1_n_600);
  L1_g29018 : OAI211D1BWP7T port map(A1 => L1_n_536, A2 => L1_n_557, B => L1_n_563, C => L1_n_537, ZN => L1_n_603);
  L1_g29019 : OAI21D0BWP7T port map(A1 => L1_n_551, A2 => L1_n_547, B => L1_n_580, ZN => L1_n_599);
  L1_g29020 : ND2D1BWP7T port map(A1 => L1_n_587, A2 => L1_n_485, ZN => L1_n_602);
  L1_g29021 : ND2D1BWP7T port map(A1 => L1_n_587, A2 => L1_n_534, ZN => L1_n_601);
  L1_g29022 : INVD0BWP7T port map(I => L1_n_596, ZN => L1_n_597);
  L1_g29023 : OAI22D0BWP7T port map(A1 => L1_n_567, A2 => L1_n_498, B1 => L1_n_549, B2 => L1_n_500, ZN => L1_n_594);
  L1_g29025 : AO21D0BWP7T port map(A1 => L1_n_550, A2 => L1_n_528, B => L1_n_577, Z => L1_n_592);
  L1_g29026 : AOI21D0BWP7T port map(A1 => L1_n_565, A2 => L1_n_489, B => L1_n_589, ZN => L1_n_598);
  L1_g29027 : AOI211D1BWP7T port map(A1 => L1_n_560, A2 => L1_n_486, B => L1_n_568, C => L1_n_71, ZN => L1_n_596);
  L1_g29028 : OAI21D0BWP7T port map(A1 => L1_n_571, A2 => L1_n_489, B => L1_n_588, ZN => L1_n_595);
  L1_g29029 : IND4D0BWP7T port map(A1 => L1_n_536, B1 => L1_n_519, B2 => L1_n_516, B3 => L1_n_540, ZN => L1_n_586);
  L1_g29030 : AOI221D0BWP7T port map(A1 => L1_n_549, A2 => L1_n_500, B1 => L1_n_490, B2 => L1_range_state_out(0), C => L1_n_533, ZN => L1_n_585);
  L1_g29031 : OA221D0BWP7T port map(A1 => L1_n_542, A2 => L1_n_65, B1 => L1_n_64, B2 => L1_n_504, C => L1_n_543, Z => L1_n_584);
  L1_g29032 : NR2XD0BWP7T port map(A1 => L1_n_566, A2 => L1_n_531, ZN => L1_n_583);
  L1_g29033 : AOI221D0BWP7T port map(A1 => L1_n_546, A2 => L1_n_64, B1 => L1_n_494, B2 => L1_n_65, C => L1_n_544, ZN => L1_n_591);
  L1_g29035 : NR2D1BWP7T port map(A1 => L1_n_565, A2 => L1_n_489, ZN => L1_n_589);
  L1_g29036 : ND2D1BWP7T port map(A1 => L1_n_571, A2 => L1_n_489, ZN => L1_n_588);
  L1_g29037 : ND2D1BWP7T port map(A1 => L1_n_569, A2 => L1_n_64, ZN => L1_n_587);
  L1_g29038 : OAI31D0BWP7T port map(A1 => L1_n_548, A2 => L1_n_538, A3 => L1_n_539, B => L1_n_528, ZN => L1_n_580);
  L1_g29039 : AO21D0BWP7T port map(A1 => L1_n_561, A2 => L1_n_487, B => L1_n_564, Z => L1_n_579);
  L1_g29040 : OR4D1BWP7T port map(A1 => L1_n_519, A2 => L1_n_488, A3 => L1_n_543, A4 => L1_n_537, Z => L1_n_578);
  L1_g29041 : AOI21D0BWP7T port map(A1 => L1_n_515, A2 => L1_n_65, B => L1_n_562, ZN => L1_n_577);
  L1_g29042 : MAOI22D0BWP7T port map(A1 => L1_n_556, A2 => L1_n_542, B1 => L1_n_504, B2 => L1_n_38, ZN => L1_n_576);
  L1_g29043 : AO211D0BWP7T port map(A1 => L1_n_487, A2 => L1_n_499, B => L1_n_558, C => L1_n_531, Z => L1_n_575);
  L1_g29044 : MOAI22D0BWP7T port map(A1 => L1_n_557, A2 => L1_n_508, B1 => L1_n_557, B2 => L1_n_508, ZN => L1_n_582);
  L1_g29046 : MAOI222D1BWP7T port map(A => L1_n_555, B => L1_n_541, C => L1_n_501, ZN => L1_n_573);
  L1_g29047 : AOI31D0BWP7T port map(A1 => L1_n_545, A2 => L1_n_530, A3 => L1_n_486, B => L1_range_state_out(0), ZN => L1_n_581);
  L1_g29048 : NR2XD0BWP7T port map(A1 => L1_n_560, A2 => L1_n_486, ZN => L1_n_568);
  L1_g29050 : OR2D1BWP7T port map(A1 => L1_n_559, A2 => L1_n_65, Z => L1_n_571);
  L1_g29051 : ND2D1BWP7T port map(A1 => L1_n_552, A2 => L1_n_508, ZN => L1_n_570);
  L1_g29052 : ND2D1BWP7T port map(A1 => L1_n_558, A2 => L1_n_531, ZN => L1_n_569);
  L1_g29053 : ND2D1BWP7T port map(A1 => L1_n_557, A2 => L1_n_518, ZN => L1_n_563);
  L1_g29054 : OAI22D0BWP7T port map(A1 => L1_n_550, A2 => L1_n_528, B1 => L1_n_515, B2 => L1_n_65, ZN => L1_n_562);
  L1_g29055 : MOAI22D0BWP7T port map(A1 => L1_n_533, A2 => L1_n_494, B1 => L1_n_533, B2 => L1_n_494, ZN => L1_n_567);
  L1_g29056 : ND2D1BWP7T port map(A1 => L1_n_558, A2 => L1_n_64, ZN => L1_n_566);
  L1_g29057 : AOI21D0BWP7T port map(A1 => L1_n_535, A2 => L1_n_543, B => L1_range_state_out(0), ZN => L1_n_565);
  L1_g29058 : NR2D1BWP7T port map(A1 => L1_n_561, A2 => L1_n_487, ZN => L1_n_564);
  L1_g29059 : INVD0BWP7T port map(I => L1_n_557, ZN => L1_n_556);
  L1_g29060 : ND2D1BWP7T port map(A1 => L1_n_545, A2 => L1_n_38, ZN => L1_n_561);
  L1_g29061 : NR2D1BWP7T port map(A1 => L1_n_546, A2 => L1_n_65, ZN => L1_n_560);
  L1_g29062 : INR2XD0BWP7T port map(A1 => L1_n_542, B1 => L1_n_537, ZN => L1_n_559);
  L1_g29063 : NR2D1BWP7T port map(A1 => L1_n_546, A2 => L1_n_486, ZN => L1_n_558);
  L1_g29064 : ND2D1BWP7T port map(A1 => L1_n_543, A2 => L1_n_38, ZN => L1_n_557);
  L1_g29065 : NR2D0BWP7T port map(A1 => L1_n_539, A2 => L1_n_538, ZN => L1_n_551);
  L1_g29066 : MAOI22D0BWP7T port map(A1 => L1_n_490, A2 => L1_n_65, B1 => L1_n_490, B2 => L1_n_65, ZN => L1_n_555);
  L1_g29067 : ND3D0BWP7T port map(A1 => L1_n_513, A2 => L1_n_510, A3 => L1_n_489, ZN => L1_n_554);
  L1_g29068 : ND2D1BWP7T port map(A1 => L1_n_534, A2 => L1_n_512, ZN => L1_n_553);
  L1_g29069 : AN2D1BWP7T port map(A1 => L1_n_542, A2 => L1_n_64, Z => L1_n_552);
  L1_g29070 : CKND1BWP7T port map(I => L1_n_547, ZN => L1_n_548);
  L1_g29071 : INVD0BWP7T port map(I => L1_n_545, ZN => L1_n_544);
  L1_g29072 : AN2D0BWP7T port map(A1 => L1_n_519, A2 => L1_n_529, Z => L1_n_550);
  L1_g29073 : IND2D1BWP7T port map(A1 => L1_n_506, B1 => L1_n_499, ZN => L1_n_549);
  L1_g29074 : IND2D1BWP7T port map(A1 => L1_n_499, B1 => L1_n_506, ZN => L1_n_541);
  L1_g29075 : NR2XD0BWP7T port map(A1 => L1_n_519, A2 => L1_n_529, ZN => L1_n_547);
  L1_g29076 : NR2XD0BWP7T port map(A1 => L1_n_494, A2 => L1_n_491, ZN => L1_n_546);
  L1_g29077 : ND2D1BWP7T port map(A1 => L1_n_494, A2 => L1_n_491, ZN => L1_n_545);
  L1_g29078 : IND2D1BWP7T port map(A1 => L1_n_504, B1 => L1_n_515, ZN => L1_n_543);
  L1_g29079 : IND2D1BWP7T port map(A1 => L1_n_515, B1 => L1_n_504, ZN => L1_n_542);
  L1_g29080 : INVD0BWP7T port map(I => L1_n_535, ZN => L1_n_536);
  L1_g29081 : INVD0BWP7T port map(I => L1_n_531, ZN => L1_n_530);
  L1_g29082 : NR2XD0BWP7T port map(A1 => L1_n_513, A2 => L1_n_510, ZN => L1_n_540);
  L1_g29083 : NR2XD0BWP7T port map(A1 => L1_n_515, A2 => L1_n_38, ZN => L1_n_539);
  L1_g29084 : CKAN2D1BWP7T port map(A1 => L1_n_515, A2 => L1_n_38, Z => L1_n_538);
  L1_g29085 : ND2D1BWP7T port map(A1 => L1_n_508, A2 => L1_n_518, ZN => L1_n_537);
  L1_g29086 : NR2D1BWP7T port map(A1 => L1_n_508, A2 => L1_n_518, ZN => L1_n_535);
  L1_g29087 : INR2D1BWP7T port map(A1 => L1_n_514, B1 => L1_n_484, ZN => L1_n_534);
  L1_g29088 : NR2XD0BWP7T port map(A1 => L1_n_490, A2 => L1_range_state_out(0), ZN => L1_n_533);
  L1_g29089 : ND3D0BWP7T port map(A1 => L1_n_482, A2 => L1_n_281, A3 => L1_n_215, ZN => L1_n_532);
  L1_g29090 : ND3D0BWP7T port map(A1 => L1_n_483, A2 => L1_n_190, A3 => L1_n_187, ZN => L1_n_531);
  L1_g29091 : INVD1BWP7T port map(I => L1_n_525, ZN => L1_n_524);
  L1_g29092 : INVD0BWP7T port map(I => L1_n_517, ZN => L1_n_516);
  L1_g29093 : INVD1BWP7T port map(I => L1_n_512, ZN => L1_n_511);
  L1_g29094 : INVD1BWP7T port map(I => L1_n_510, ZN => L1_n_509);
  L1_g29096 : ND3D0BWP7T port map(A1 => L1_n_465, A2 => L1_n_240, A3 => L1_n_161, ZN => L1_n_529);
  L1_g29097 : ND3D0BWP7T port map(A1 => L1_n_459, A2 => L1_n_246, A3 => L1_n_245, ZN => L1_n_528);
  L1_g29098 : ND3D0BWP7T port map(A1 => L1_n_472, A2 => L1_n_267, A3 => L1_n_265, ZN => L1_n_527);
  L1_g29099 : ND3D0BWP7T port map(A1 => L1_n_476, A2 => L1_n_294, A3 => L1_n_295, ZN => L1_n_526);
  L1_g29100 : ND3D0BWP7T port map(A1 => L1_n_478, A2 => L1_n_302, A3 => L1_n_304, ZN => L1_n_525);
  L1_g29101 : ND3D0BWP7T port map(A1 => L1_n_467, A2 => L1_n_252, A3 => L1_n_251, ZN => L1_n_523);
  L1_g29102 : ND3D0BWP7T port map(A1 => L1_n_481, A2 => L1_n_279, A3 => L1_n_317, ZN => L1_n_522);
  L1_g29103 : AN3D1BWP7T port map(A1 => L1_n_469, A2 => L1_n_259, A3 => L1_n_260, Z => L1_n_521);
  L1_g29104 : ND3D0BWP7T port map(A1 => L1_n_473, A2 => L1_n_272, A3 => L1_n_271, ZN => L1_n_520);
  L1_g29105 : AN3D1BWP7T port map(A1 => L1_n_479, A2 => L1_n_303, A3 => L1_n_301, Z => L1_n_519);
  L1_g29106 : ND3D0BWP7T port map(A1 => L1_n_475, A2 => L1_n_276, A3 => L1_n_280, ZN => L1_n_518);
  L1_g29107 : ND3D0BWP7T port map(A1 => L1_n_477, A2 => L1_n_293, A3 => L1_n_292, ZN => L1_n_517);
  L1_g29108 : ND3D0BWP7T port map(A1 => L1_n_480, A2 => L1_n_310, A3 => L1_n_309, ZN => L1_n_515);
  L1_g29109 : ND3D0BWP7T port map(A1 => L1_n_463, A2 => L1_n_224, A3 => L1_n_222, ZN => L1_n_514);
  L1_g29110 : ND3D0BWP7T port map(A1 => L1_n_470, A2 => L1_n_257, A3 => L1_n_258, ZN => L1_n_513);
  L1_g29111 : ND3D0BWP7T port map(A1 => L1_n_464, A2 => L1_n_235, A3 => L1_n_234, ZN => L1_n_512);
  L1_g29112 : ND3D0BWP7T port map(A1 => L1_n_468, A2 => L1_n_247, A3 => L1_n_248, ZN => L1_n_510);
  L1_g29113 : ND3D0BWP7T port map(A1 => L1_n_471, A2 => L1_n_266, A3 => L1_n_268, ZN => L1_n_508);
  L1_g29114 : INVD0BWP7T port map(I => L1_n_500, ZN => L1_n_501);
  L1_g29115 : INVD0BWP7T port map(I => L1_n_496, ZN => L1_n_495);
  L1_g29116 : INVD1BWP7T port map(I => L1_n_492, ZN => L1_n_493);
  L1_g29117 : INVD1BWP7T port map(I => L1_n_491, ZN => L1_n_490);
  L1_g29118 : INVD0BWP7T port map(I => L1_n_489, ZN => L1_n_488);
  L1_g29119 : INVD1BWP7T port map(I => L1_n_487, ZN => L1_n_486);
  L1_g29120 : INVD1BWP7T port map(I => L1_n_485, ZN => L1_n_484);
  L1_g29121 : AOI221D0BWP7T port map(A1 => L1_n_101, A2 => y_4(4), B1 => L1_n_83, B2 => y_12(4), C => L1_n_446, ZN => L1_n_483);
  L1_g29122 : AOI221D0BWP7T port map(A1 => L1_n_101, A2 => y_4(8), B1 => L1_n_86, B2 => y_14(8), C => L1_n_447, ZN => L1_n_482);
  L1_g29123 : ND3D0BWP7T port map(A1 => L1_n_457, A2 => L1_n_189, A3 => L1_n_188, ZN => L1_n_506);
  L1_g29124 : AN3D1BWP7T port map(A1 => L1_n_466, A2 => L1_n_209, A3 => L1_n_210, Z => L1_n_505);
  L1_g29125 : AN3D1BWP7T port map(A1 => L1_n_452, A2 => L1_n_165, A3 => L1_n_169, Z => L1_n_504);
  L1_g29126 : ND3D0BWP7T port map(A1 => L1_n_461, A2 => L1_n_221, A3 => L1_n_205, ZN => L1_n_503);
  L1_g29127 : ND3D0BWP7T port map(A1 => L1_n_460, A2 => L1_n_216, A3 => L1_n_217, ZN => L1_n_502);
  L1_g29128 : ND4D0BWP7T port map(A1 => L1_n_448, A2 => L1_n_195, A3 => L1_n_196, A4 => L1_n_307, ZN => L1_n_500);
  L1_g29129 : ND3D0BWP7T port map(A1 => L1_n_455, A2 => L1_n_175, A3 => L1_n_179, ZN => L1_n_499);
  L1_g29130 : ND4D0BWP7T port map(A1 => L1_n_449, A2 => L1_n_202, A3 => L1_n_203, A4 => L1_n_172, ZN => L1_n_498);
  L1_g29131 : ND4D0BWP7T port map(A1 => L1_n_450, A2 => L1_n_166, A3 => L1_n_230, A4 => L1_n_231, ZN => L1_n_497);
  L1_g29132 : ND4D0BWP7T port map(A1 => L1_n_451, A2 => L1_n_287, A3 => L1_n_286, A4 => L1_n_284, ZN => L1_n_496);
  L1_g29133 : ND3D0BWP7T port map(A1 => L1_n_453, A2 => L1_n_168, A3 => L1_n_167, ZN => L1_n_494);
  L1_g29134 : ND3D0BWP7T port map(A1 => L1_n_462, A2 => L1_n_225, A3 => L1_n_226, ZN => L1_n_492);
  L1_g29135 : ND3D0BWP7T port map(A1 => L1_n_474, A2 => L1_n_314, A3 => L1_n_313, ZN => L1_n_491);
  L1_g29136 : ND3D0BWP7T port map(A1 => L1_n_454, A2 => L1_n_184, A3 => L1_n_191, ZN => L1_n_489);
  L1_g29137 : ND3D0BWP7T port map(A1 => L1_n_456, A2 => L1_n_178, A3 => L1_n_177, ZN => L1_n_487);
  L1_g29138 : ND3D0BWP7T port map(A1 => L1_n_458, A2 => L1_n_233, A3 => L1_n_201, ZN => L1_n_485);
  L1_g29139 : AOI221D0BWP7T port map(A1 => L1_n_107, A2 => x_11(7), B1 => L1_n_108, B2 => x_7(7), C => L1_n_437, ZN => L1_n_481);
  L1_g29140 : AOI221D0BWP7T port map(A1 => L1_n_103, A2 => x_6(1), B1 => L1_n_82, B2 => x_8(1), C => L1_n_442, ZN => L1_n_480);
  L1_g29141 : AOI221D0BWP7T port map(A1 => L1_n_101, A2 => x_4(0), B1 => L1_n_83, B2 => x_12(0), C => L1_n_440, ZN => L1_n_479);
  L1_g29142 : AOI221D0BWP7T port map(A1 => L1_n_85, A2 => x_2(8), B1 => L1_n_102, B2 => x_14(8), C => L1_n_445, ZN => L1_n_478);
  L1_g29143 : AOI221D0BWP7T port map(A1 => L1_n_82, A2 => x_8(8), B1 => L1_n_103, B2 => x_6(8), C => L1_n_438, ZN => L1_n_477);
  L1_g29144 : AOI221D0BWP7T port map(A1 => L1_n_109, A2 => y_8(8), B1 => L1_n_111, B2 => y_0(8), C => L1_n_439, ZN => L1_n_476);
  L1_g29145 : AOI221D0BWP7T port map(A1 => L1_n_101, A2 => x_4(4), B1 => L1_n_86, B2 => x_14(4), C => L1_n_435, ZN => L1_n_475);
  L1_g29146 : AOI221D0BWP7T port map(A1 => L1_n_88, A2 => y_1(1), B1 => L1_n_91, B2 => y_7(1), C => L1_n_443, ZN => L1_n_474);
  L1_g29147 : AOI221D0BWP7T port map(A1 => L1_n_109, A2 => x_8(5), B1 => L1_n_111, B2 => x_0(5), C => L1_n_436, ZN => L1_n_473);
  L1_g29148 : AOI221D0BWP7T port map(A1 => L1_n_107, A2 => x_11(4), B1 => L1_n_108, B2 => x_7(4), C => L1_n_434, ZN => L1_n_472);
  L1_g29149 : AOI221D0BWP7T port map(A1 => L1_n_101, A2 => x_4(3), B1 => L1_n_86, B2 => x_14(3), C => L1_n_433, ZN => L1_n_471);
  L1_g29150 : AOI221D0BWP7T port map(A1 => L1_n_101, A2 => x_4(7), B1 => L1_n_86, B2 => x_14(7), C => L1_n_431, ZN => L1_n_470);
  L1_g29151 : AOI221D0BWP7T port map(A1 => L1_n_109, A2 => x_8(3), B1 => L1_n_111, B2 => x_0(3), C => L1_n_432, ZN => L1_n_469);
  L1_g29152 : AOI221D0BWP7T port map(A1 => L1_n_101, A2 => x_4(6), B1 => L1_n_86, B2 => x_14(6), C => L1_n_428, ZN => L1_n_468);
  L1_g29153 : AOI221D0BWP7T port map(A1 => L1_n_85, A2 => x_2(2), B1 => L1_n_99, B2 => x_15(2), C => L1_n_430, ZN => L1_n_467);
  L1_g29154 : AOI221D0BWP7T port map(A1 => L1_n_85, A2 => y_2(3), B1 => L1_n_99, B2 => y_15(3), C => L1_n_420, ZN => L1_n_466);
  L1_g29155 : AOI221D0BWP7T port map(A1 => L1_n_105, A2 => x_12(0), B1 => L1_n_112, B2 => x_4(0), C => L1_n_427, ZN => L1_n_465);
  L1_g29156 : AOI221D0BWP7T port map(A1 => L1_n_101, A2 => y_4(7), B1 => L1_n_83, B2 => y_12(7), C => L1_n_426, ZN => L1_n_464);
  L1_g29157 : AOI221D0BWP7T port map(A1 => L1_n_101, A2 => y_4(6), B1 => L1_n_92, B2 => y_3(6), C => L1_n_424, ZN => L1_n_463);
  L1_g29158 : AOI221D0BWP7T port map(A1 => L1_n_81, A2 => y_10(7), B1 => L1_n_108, B2 => y_7(7), C => L1_n_425, ZN => L1_n_462);
  L1_g29159 : AOI221D0BWP7T port map(A1 => L1_n_109, A2 => y_8(5), B1 => L1_n_111, B2 => y_0(5), C => L1_n_423, ZN => L1_n_461);
  L1_g29160 : AOI221D0BWP7T port map(A1 => L1_n_102, A2 => y_14(4), B1 => L1_n_111, B2 => y_0(4), C => L1_n_422, ZN => L1_n_460);
  L1_g29161 : AOI221D0BWP7T port map(A1 => L1_n_107, A2 => x_11(1), B1 => L1_n_108, B2 => x_7(1), C => L1_n_429, ZN => L1_n_459);
  L1_g29162 : AOI221D0BWP7T port map(A1 => L1_n_101, A2 => y_4(5), B1 => L1_n_92, B2 => y_3(5), C => L1_n_419, ZN => L1_n_458);
  L1_g29163 : AOI221D0BWP7T port map(A1 => L1_n_106, A2 => y_3(0), B1 => L1_n_102, B2 => y_14(0), C => L1_n_418, ZN => L1_n_457);
  L1_g29164 : AOI221D0BWP7T port map(A1 => L1_n_101, A2 => y_4(3), B1 => L1_n_83, B2 => y_12(3), C => L1_n_417, ZN => L1_n_456);
  L1_g29165 : AOI221D0BWP7T port map(A1 => L1_n_103, A2 => y_6(0), B1 => L1_n_88, B2 => y_1(0), C => L1_n_416, ZN => L1_n_455);
  L1_g29166 : AOI221D0BWP7T port map(A1 => L1_n_101, A2 => x_4(5), B1 => L1_n_113, B2 => x_15(5), C => L1_n_421, ZN => L1_n_454);
  L1_g29167 : AOI221D0BWP7T port map(A1 => L1_n_113, A2 => y_15(2), B1 => L1_n_101, B2 => y_4(2), C => L1_n_415, ZN => L1_n_453);
  L1_g29168 : AOI221D0BWP7T port map(A1 => L1_n_101, A2 => x_4(2), B1 => L1_n_94, B2 => x_13(2), C => L1_n_414, ZN => L1_n_452);
  L1_g29169 : AOI221D0BWP7T port map(A1 => L1_n_96, A2 => x_5(6), B1 => L1_n_110, B2 => x_13(6), C => L1_n_441, ZN => L1_n_451);
  L1_g29170 : AOI221D0BWP7T port map(A1 => L1_n_81, A2 => y_10(6), B1 => L1_n_84, B2 => y_6(6), C => L1_n_444, ZN => L1_n_450);
  L1_g29171 : AOI221D0BWP7T port map(A1 => L1_n_85, A2 => y_2(2), B1 => L1_n_99, B2 => y_15(2), C => L1_n_395, ZN => L1_n_449);
  L1_g29172 : AOI221D0BWP7T port map(A1 => L1_n_85, A2 => y_2(1), B1 => L1_n_99, B2 => y_15(1), C => L1_n_394, ZN => L1_n_448);
  L1_g29173 : ND4D0BWP7T port map(A1 => L1_n_405, A2 => L1_n_212, A3 => L1_n_211, A4 => L1_n_208, ZN => L1_n_447);
  L1_g29174 : ND4D0BWP7T port map(A1 => L1_n_404, A2 => L1_n_182, A3 => L1_n_183, A4 => L1_n_180, ZN => L1_n_446);
  L1_g29175 : ND4D0BWP7T port map(A1 => L1_n_344, A2 => L1_n_376, A3 => L1_n_300, A4 => L1_n_298, ZN => L1_n_445);
  L1_g29176 : ND4D0BWP7T port map(A1 => L1_n_360, A2 => L1_n_227, A3 => L1_n_228, A4 => L1_n_152, ZN => L1_n_444);
  L1_g29177 : ND4D0BWP7T port map(A1 => L1_n_346, A2 => L1_n_378, A3 => L1_n_312, A4 => L1_n_311, ZN => L1_n_443);
  L1_g29178 : ND4D0BWP7T port map(A1 => L1_n_377, A2 => L1_n_345, A3 => L1_n_305, A4 => L1_n_306, ZN => L1_n_442);
  L1_g29179 : ND4D0BWP7T port map(A1 => L1_n_372, A2 => L1_n_283, A3 => L1_n_282, A4 => L1_n_150, ZN => L1_n_441);
  L1_g29180 : ND4D0BWP7T port map(A1 => L1_n_299, A2 => L1_n_296, A3 => L1_n_375, A4 => L1_n_343, ZN => L1_n_440);
  L1_g29181 : ND4D0BWP7T port map(A1 => L1_n_342, A2 => L1_n_374, A3 => L1_n_290, A4 => L1_n_291, ZN => L1_n_439);
  L1_g29182 : ND4D0BWP7T port map(A1 => L1_n_289, A2 => L1_n_285, A3 => L1_n_373, A4 => L1_n_341, ZN => L1_n_438);
  L1_g29199 : ND4D0BWP7T port map(A1 => L1_n_340, A2 => L1_n_371, A3 => L1_n_277, A4 => L1_n_275, ZN => L1_n_437);
  L1_g29200 : ND4D0BWP7T port map(A1 => L1_n_338, A2 => L1_n_369, A3 => L1_n_269, A4 => L1_n_270, ZN => L1_n_436);
  L1_g29201 : ND4D0BWP7T port map(A1 => L1_n_339, A2 => L1_n_370, A3 => L1_n_273, A4 => L1_n_274, ZN => L1_n_435);
  L1_g29202 : ND4D0BWP7T port map(A1 => L1_n_337, A2 => L1_n_368, A3 => L1_n_262, A4 => L1_n_263, ZN => L1_n_434);
  L1_g29203 : ND4D0BWP7T port map(A1 => L1_n_367, A2 => L1_n_336, A3 => L1_n_261, A4 => L1_n_264, ZN => L1_n_433);
  L1_g29204 : ND4D0BWP7T port map(A1 => L1_n_335, A2 => L1_n_366, A3 => L1_n_255, A4 => L1_n_256, ZN => L1_n_432);
  L1_g29205 : ND4D0BWP7T port map(A1 => L1_n_364, A2 => L1_n_334, A3 => L1_n_254, A4 => L1_n_253, ZN => L1_n_431);
  L1_g29206 : ND4D0BWP7T port map(A1 => L1_n_333, A2 => L1_n_365, A3 => L1_n_250, A4 => L1_n_249, ZN => L1_n_430);
  L1_g29207 : ND4D0BWP7T port map(A1 => L1_n_332, A2 => L1_n_363, A3 => L1_n_244, A4 => L1_n_243, ZN => L1_n_429);
  L1_g29208 : ND4D0BWP7T port map(A1 => L1_n_362, A2 => L1_n_331, A3 => L1_n_242, A4 => L1_n_241, ZN => L1_n_428);
  L1_g29209 : ND4D0BWP7T port map(A1 => L1_n_330, A2 => L1_n_361, A3 => L1_n_237, A4 => L1_n_236, ZN => L1_n_427);
  L1_g29210 : ND4D0BWP7T port map(A1 => L1_n_232, A2 => L1_n_229, A3 => L1_n_329, A4 => L1_n_359, ZN => L1_n_426);
  L1_g29211 : ND4D0BWP7T port map(A1 => L1_n_328, A2 => L1_n_358, A3 => L1_n_238, A4 => L1_n_223, ZN => L1_n_425);
  L1_g29212 : ND4D0BWP7T port map(A1 => L1_n_356, A2 => L1_n_327, A3 => L1_n_219, A4 => L1_n_220, ZN => L1_n_424);
  L1_g29213 : ND4D0BWP7T port map(A1 => L1_n_326, A2 => L1_n_357, A3 => L1_n_218, A4 => L1_n_204, ZN => L1_n_423);
  L1_g29214 : ND4D0BWP7T port map(A1 => L1_n_325, A2 => L1_n_355, A3 => L1_n_214, A4 => L1_n_213, ZN => L1_n_422);
  L1_g29215 : ND4D0BWP7T port map(A1 => L1_n_349, A2 => L1_n_320, A3 => L1_n_288, A4 => L1_n_176, ZN => L1_n_421);
  L1_g29216 : ND4D0BWP7T port map(A1 => L1_n_324, A2 => L1_n_354, A3 => L1_n_206, A4 => L1_n_207, ZN => L1_n_420);
  L1_g29217 : ND4D0BWP7T port map(A1 => L1_n_353, A2 => L1_n_323, A3 => L1_n_197, A4 => L1_n_308, ZN => L1_n_419);
  L1_g29218 : ND4D0BWP7T port map(A1 => L1_n_322, A2 => L1_n_352, A3 => L1_n_186, A4 => L1_n_185, ZN => L1_n_418);
  L1_g29219 : ND4D0BWP7T port map(A1 => L1_n_321, A2 => L1_n_351, A3 => L1_n_174, A4 => L1_n_173, ZN => L1_n_417);
  L1_g29220 : ND4D0BWP7T port map(A1 => L1_n_350, A2 => L1_n_319, A3 => L1_n_170, A4 => L1_n_171, ZN => L1_n_416);
  L1_g29221 : ND4D0BWP7T port map(A1 => L1_n_318, A2 => L1_n_348, A3 => L1_n_164, A4 => L1_n_163, ZN => L1_n_415);
  L1_g29222 : ND4D0BWP7T port map(A1 => L1_n_347, A2 => L1_n_379, A3 => L1_n_162, A4 => L1_n_239, ZN => L1_n_414);
  L1_g29223 : IOA21D1BWP7T port map(A1 => L1_n_158, A2 => L1_n_46, B => L1_n_389, ZN => L1_n_413);
  L1_g29224 : IOA21D1BWP7T port map(A1 => L1_n_0, A2 => L1_n_46, B => L1_n_385, ZN => L1_n_412);
  L1_g29225 : MOAI22D0BWP7T port map(A1 => L1_n_157, A2 => L1_n_702, B1 => L1_n_316, B2 => FE_PHN9_L1_n_25, ZN => L1_n_411);
  L1_g29226 : IOA21D1BWP7T port map(A1 => L1_n_156, A2 => L1_n_46, B => L1_n_384, ZN => L1_n_410);
  L1_g29227 : IOA21D1BWP7T port map(A1 => L1_n_158, A2 => L1_n_68, B => L1_n_388, ZN => L1_n_409);
  L1_g29228 : IOA21D1BWP7T port map(A1 => L1_n_0, A2 => L1_n_68, B => L1_n_382, ZN => L1_n_408);
  L1_g29229 : IOA21D1BWP7T port map(A1 => L1_n_156, A2 => L1_n_68, B => L1_n_381, ZN => L1_n_407);
  L1_g29230 : IOA21D1BWP7T port map(A1 => L1_n_156, A2 => L1_n_60, B => L1_n_391, ZN => L1_n_406);
  L1_g29231 : AOI222D0BWP7T port map(A1 => L1_n_147, A2 => L1_n_46, B1 => L1_n_94, B2 => y_13(8), C1 => L1_n_113, C2 => y_15(8), ZN => L1_n_405);
  L1_g29232 : AOI222D0BWP7T port map(A1 => L1_n_151, A2 => L1_n_46, B1 => L1_n_94, B2 => y_13(4), C1 => L1_n_113, C2 => y_15(4), ZN => L1_n_404);
  L1_g29233 : IOA21D1BWP7T port map(A1 => L1_n_158, A2 => L1_n_60, B => L1_n_392, ZN => L1_n_403);
  L1_g29234 : IOA21D1BWP7T port map(A1 => L1_n_0, A2 => L1_n_60, B => L1_n_380, ZN => L1_n_402);
  L1_g29235 : IOA21D1BWP7T port map(A1 => L1_n_0, A2 => L1_n_41, B => L1_n_386, ZN => L1_n_401);
  L1_g29236 : OAI21D0BWP7T port map(A1 => L1_n_159, A2 => L1_n_702, B => L1_n_393, ZN => L1_n_400);
  L1_g29237 : OAI21D0BWP7T port map(A1 => L1_n_159, A2 => L1_n_47, B => L1_n_387, ZN => L1_n_399);
  L1_g29238 : AO22D0BWP7T port map(A1 => L1_n_278, A2 => FE_PHN4_L1_n_21, B1 => L1_n_41, B2 => L1_n_158, Z => L1_n_398);
  L1_g29239 : OAI21D0BWP7T port map(A1 => L1_n_159, A2 => L1_n_69, B => L1_n_383, ZN => L1_n_397);
  L1_g29240 : OAI21D0BWP7T port map(A1 => L1_n_159, A2 => L1_n_61, B => L1_n_390, ZN => L1_n_396);
  L1_g29241 : ND4D0BWP7T port map(A1 => L1_n_200, A2 => L1_n_199, A3 => L1_n_297, A4 => L1_n_198, ZN => L1_n_395);
  L1_g29242 : ND4D0BWP7T port map(A1 => L1_n_181, A2 => L1_n_193, A3 => L1_n_192, A4 => L1_n_194, ZN => L1_n_394);
  L1_g29243 : OAI21D0BWP7T port map(A1 => L1_n_1, A2 => L1_n_59, B => FE_PHN8_L1_n_19, ZN => L1_n_393);
  L1_g29244 : OAI21D0BWP7T port map(A1 => L1_n_115, A2 => L1_n_154, B => FE_PHN6_L1_n_30, ZN => L1_n_392);
  L1_g29245 : OAI21D0BWP7T port map(A1 => L1_n_115, A2 => L1_n_155, B => FE_PHN3_L1_n_34, ZN => L1_n_391);
  L1_g29246 : OAI21D0BWP7T port map(A1 => L1_n_115, A2 => L1_n_1, B => FE_PHN12_L1_n_28, ZN => L1_n_390);
  L1_g29247 : OAI21D0BWP7T port map(A1 => L1_n_114, A2 => L1_n_154, B => FE_PHN13_L1_n_22, ZN => L1_n_389);
  L1_g29248 : OAI21D0BWP7T port map(A1 => L1_n_154, A2 => L1_n_116, B => FE_PHN5_L1_n_29, ZN => L1_n_388);
  L1_g29249 : OAI21D0BWP7T port map(A1 => L1_n_114, A2 => L1_n_1, B => FE_PHN10_L1_n_20, ZN => L1_n_387);
  L1_g29250 : OAI21D0BWP7T port map(A1 => L1_n_160, A2 => L1_n_59, B => FE_PHN16_L1_n_23, ZN => L1_n_386);
  L1_g29251 : OAI21D0BWP7T port map(A1 => L1_n_114, A2 => L1_n_160, B => FE_PHN14_L1_n_24, ZN => L1_n_385);
  L1_g29252 : OAI21D0BWP7T port map(A1 => L1_n_114, A2 => L1_n_155, B => FE_PHN1_L1_n_26, ZN => L1_n_384);
  L1_g29253 : OAI21D0BWP7T port map(A1 => L1_n_1, A2 => L1_n_116, B => FE_PHN11_L1_n_27, ZN => L1_n_383);
  L1_g29254 : OAI21D0BWP7T port map(A1 => L1_n_116, A2 => L1_n_160, B => FE_PHN7_L1_n_31, ZN => L1_n_382);
  L1_g29255 : OAI21D0BWP7T port map(A1 => L1_n_116, A2 => L1_n_155, B => L1_n_33, ZN => L1_n_381);
  L1_g29256 : OAI21D0BWP7T port map(A1 => L1_n_115, A2 => L1_n_160, B => FE_PHN2_L1_n_32, ZN => L1_n_380);
  L1_g29257 : AOI222D0BWP7T port map(A1 => L1_n_104, A2 => x_2(2), B1 => L1_n_87, B2 => x_10(2), C1 => L1_n_86, C2 => x_14(2), ZN => L1_n_379);
  L1_g29258 : AOI222D0BWP7T port map(A1 => L1_n_104, A2 => y_2(1), B1 => L1_n_87, B2 => y_10(1), C1 => L1_n_86, C2 => y_14(1), ZN => L1_n_378);
  L1_g29259 : AOI222D0BWP7T port map(A1 => L1_n_104, A2 => x_2(1), B1 => L1_n_92, B2 => x_3(1), C1 => L1_n_94, C2 => x_13(1), ZN => L1_n_377);
  L1_g29260 : AOI222D0BWP7T port map(A1 => L1_n_109, A2 => x_8(8), B1 => L1_n_105, B2 => x_12(8), C1 => L1_n_84, C2 => x_6(8), ZN => L1_n_376);
  L1_g29261 : AOI222D0BWP7T port map(A1 => L1_n_104, A2 => x_2(0), B1 => L1_n_97, B2 => x_11(0), C1 => L1_n_113, C2 => x_15(0), ZN => L1_n_375);
  L1_g29262 : AOI222D0BWP7T port map(A1 => L1_n_107, A2 => y_11(8), B1 => L1_n_99, B2 => y_15(8), C1 => L1_n_84, C2 => y_6(8), ZN => L1_n_374);
  L1_g29263 : AOI222D0BWP7T port map(A1 => L1_n_104, A2 => x_2(8), B1 => L1_n_97, B2 => x_11(8), C1 => L1_n_113, C2 => x_15(8), ZN => L1_n_373);
  L1_g29264 : AOI222D0BWP7T port map(A1 => L1_n_85, A2 => x_2(6), B1 => L1_n_84, B2 => x_6(6), C1 => L1_n_105, C2 => x_12(6), ZN => L1_n_372);
  L1_g29265 : AOI222D0BWP7T port map(A1 => L1_n_111, A2 => x_0(7), B1 => L1_n_112, B2 => x_4(7), C1 => L1_n_84, C2 => x_6(7), ZN => L1_n_371);
  L1_g29266 : AOI222D0BWP7T port map(A1 => L1_n_104, A2 => x_2(4), B1 => L1_n_97, B2 => x_11(4), C1 => L1_n_113, C2 => x_15(4), ZN => L1_n_370);
  L1_g29267 : AOI222D0BWP7T port map(A1 => L1_n_106, A2 => x_3(5), B1 => L1_n_108, B2 => x_7(5), C1 => L1_n_84, C2 => x_6(5), ZN => L1_n_369);
  L1_g29268 : AOI222D0BWP7T port map(A1 => L1_n_111, A2 => x_0(4), B1 => L1_n_112, B2 => x_4(4), C1 => L1_n_84, C2 => x_6(4), ZN => L1_n_368);
  L1_g29269 : AOI222D0BWP7T port map(A1 => L1_n_104, A2 => x_2(3), B1 => L1_n_92, B2 => x_3(3), C1 => L1_n_94, C2 => x_13(3), ZN => L1_n_367);
  L1_g29270 : AOI222D0BWP7T port map(A1 => L1_n_107, A2 => x_11(3), B1 => L1_n_99, B2 => x_15(3), C1 => L1_n_84, C2 => x_6(3), ZN => L1_n_366);
  L1_g29271 : AOI222D0BWP7T port map(A1 => L1_n_111, A2 => x_0(2), B1 => L1_n_112, B2 => x_4(2), C1 => L1_n_84, C2 => x_6(2), ZN => L1_n_365);
  L1_g29272 : AOI222D0BWP7T port map(A1 => L1_n_104, A2 => x_2(7), B1 => L1_n_92, B2 => x_3(7), C1 => L1_n_94, C2 => x_13(7), ZN => L1_n_364);
  L1_g29273 : AOI222D0BWP7T port map(A1 => L1_n_109, A2 => x_8(1), B1 => L1_n_105, B2 => x_12(1), C1 => L1_n_84, C2 => x_6(1), ZN => L1_n_363);
  L1_g29274 : AOI222D0BWP7T port map(A1 => L1_n_104, A2 => x_2(6), B1 => L1_n_92, B2 => x_3(6), C1 => L1_n_94, C2 => x_13(6), ZN => L1_n_362);
  L1_g29275 : AOI222D0BWP7T port map(A1 => L1_n_107, A2 => x_11(0), B1 => L1_n_99, B2 => x_15(0), C1 => L1_n_84, C2 => x_6(0), ZN => L1_n_361);
  L1_g29276 : AOI222D0BWP7T port map(A1 => L1_n_95, A2 => y_1(6), B1 => L1_n_96, B2 => y_5(6), C1 => L1_n_108, C2 => y_7(6), ZN => L1_n_360);
  L1_g29277 : AOI222D0BWP7T port map(A1 => L1_n_104, A2 => y_2(7), B1 => L1_n_97, B2 => y_11(7), C1 => L1_n_113, C2 => y_15(7), ZN => L1_n_359);
  L1_g29278 : AOI222D0BWP7T port map(A1 => L1_n_111, A2 => y_0(7), B1 => L1_n_112, B2 => y_4(7), C1 => L1_n_84, C2 => y_6(7), ZN => L1_n_358);
  L1_g29279 : AOI222D0BWP7T port map(A1 => L1_n_107, A2 => y_11(5), B1 => L1_n_99, B2 => y_15(5), C1 => L1_n_84, C2 => y_6(5), ZN => L1_n_357);
  L1_g29280 : AOI222D0BWP7T port map(A1 => L1_n_104, A2 => y_2(6), B1 => L1_n_87, B2 => y_10(6), C1 => L1_n_86, C2 => y_14(6), ZN => L1_n_356);
  L1_g29281 : AOI222D0BWP7T port map(A1 => L1_n_107, A2 => y_11(4), B1 => L1_n_99, B2 => y_15(4), C1 => L1_n_84, C2 => y_6(4), ZN => L1_n_355);
  L1_g29282 : AOI222D0BWP7T port map(A1 => L1_n_111, A2 => y_0(3), B1 => L1_n_112, B2 => y_4(3), C1 => L1_n_84, C2 => y_6(3), ZN => L1_n_354);
  L1_g29283 : AOI222D0BWP7T port map(A1 => L1_n_87, A2 => y_10(5), B1 => L1_n_86, B2 => y_14(5), C1 => L1_n_104, C2 => y_2(5), ZN => L1_n_353);
  L1_g29284 : AOI222D0BWP7T port map(A1 => L1_n_111, A2 => y_0(0), B1 => L1_n_112, B2 => y_4(0), C1 => L1_n_84, C2 => y_6(0), ZN => L1_n_352);
  L1_g29285 : AOI222D0BWP7T port map(A1 => L1_n_104, A2 => y_2(3), B1 => L1_n_92, B2 => y_3(3), C1 => L1_n_94, C2 => y_13(3), ZN => L1_n_351);
  L1_g29286 : AOI222D0BWP7T port map(A1 => L1_n_104, A2 => y_2(0), B1 => L1_n_87, B2 => y_10(0), C1 => L1_n_86, C2 => y_14(0), ZN => L1_n_350);
  L1_g29287 : AOI222D0BWP7T port map(A1 => L1_n_104, A2 => x_2(5), B1 => L1_n_87, B2 => x_10(5), C1 => L1_n_86, C2 => x_14(5), ZN => L1_n_349);
  L1_g29288 : AOI222D0BWP7T port map(A1 => L1_n_104, A2 => y_2(2), B1 => L1_n_82, B2 => y_8(2), C1 => L1_n_83, C2 => y_12(2), ZN => L1_n_348);
  L1_g29289 : MAOI22D0BWP7T port map(A1 => L1_n_100, A2 => x_0(2), B1 => L1_n_143, B2 => L1_n_47, ZN => L1_n_347);
  L1_g29290 : MAOI22D0BWP7T port map(A1 => L1_n_100, A2 => y_0(1), B1 => L1_n_146, B2 => L1_n_61, ZN => L1_n_346);
  L1_g29291 : MAOI22D0BWP7T port map(A1 => L1_n_100, A2 => x_0(1), B1 => L1_n_125, B2 => L1_n_61, ZN => L1_n_345);
  L1_g29292 : MAOI22D0BWP7T port map(A1 => L1_n_106, A2 => x_3(8), B1 => L1_n_70, B2 => L1_n_129, ZN => L1_n_344);
  L1_g29293 : MAOI22D0BWP7T port map(A1 => L1_n_100, A2 => x_0(0), B1 => L1_n_139, B2 => L1_n_61, ZN => L1_n_343);
  L1_g29294 : MAOI22D0BWP7T port map(A1 => L1_n_85, A2 => y_2(8), B1 => L1_n_50, B2 => L1_n_137, ZN => L1_n_342);
  L1_g29295 : MAOI22D0BWP7T port map(A1 => L1_n_100, A2 => x_0(8), B1 => L1_n_124, B2 => L1_n_61, ZN => L1_n_341);
  L1_g29296 : MAOI22D0BWP7T port map(A1 => L1_n_106, A2 => x_3(7), B1 => L1_n_50, B2 => L1_n_133, ZN => L1_n_340);
  L1_g29297 : MAOI22D0BWP7T port map(A1 => L1_n_100, A2 => x_0(4), B1 => L1_n_132, B2 => L1_n_47, ZN => L1_n_339);
  L1_g29298 : MAOI22D0BWP7T port map(A1 => L1_n_85, A2 => x_2(5), B1 => L1_n_56, B2 => L1_n_127, ZN => L1_n_338);
  L1_g29299 : MAOI22D0BWP7T port map(A1 => L1_n_106, A2 => x_3(4), B1 => L1_n_50, B2 => L1_n_141, ZN => L1_n_337);
  L1_g29300 : MAOI22D0BWP7T port map(A1 => L1_n_100, A2 => x_0(3), B1 => L1_n_138, B2 => L1_n_61, ZN => L1_n_336);
  L1_g29301 : MAOI22D0BWP7T port map(A1 => L1_n_85, A2 => x_2(3), B1 => L1_n_56, B2 => L1_n_140, ZN => L1_n_335);
  L1_g29302 : MAOI22D0BWP7T port map(A1 => L1_n_100, A2 => x_0(7), B1 => L1_n_144, B2 => L1_n_61, ZN => L1_n_334);
  L1_g29303 : MAOI22D0BWP7T port map(A1 => L1_n_106, A2 => x_3(2), B1 => L1_n_50, B2 => L1_n_131, ZN => L1_n_333);
  L1_g29304 : MAOI22D0BWP7T port map(A1 => L1_n_106, A2 => x_3(1), B1 => L1_n_70, B2 => L1_n_123, ZN => L1_n_332);
  L1_g29305 : MAOI22D0BWP7T port map(A1 => L1_n_100, A2 => x_0(6), B1 => L1_n_130, B2 => L1_n_61, ZN => L1_n_331);
  L1_g29306 : MAOI22D0BWP7T port map(A1 => L1_n_85, A2 => x_2(0), B1 => L1_n_50, B2 => L1_n_126, ZN => L1_n_330);
  L1_g29307 : MAOI22D0BWP7T port map(A1 => L1_n_100, A2 => y_0(7), B1 => L1_n_148, B2 => L1_n_61, ZN => L1_n_329);
  L1_g29308 : MAOI22D0BWP7T port map(A1 => L1_n_85, A2 => y_2(7), B1 => L1_n_50, B2 => L1_n_128, ZN => L1_n_328);
  L1_g29309 : MAOI22D0BWP7T port map(A1 => L1_n_100, A2 => y_0(6), B1 => L1_n_122, B2 => L1_n_61, ZN => L1_n_327);
  L1_g29310 : MAOI22D0BWP7T port map(A1 => L1_n_85, A2 => y_2(5), B1 => L1_n_50, B2 => L1_n_121, ZN => L1_n_326);
  L1_g29311 : MAOI22D0BWP7T port map(A1 => L1_n_85, A2 => y_2(4), B1 => L1_n_50, B2 => L1_n_149, ZN => L1_n_325);
  L1_g29312 : MAOI22D0BWP7T port map(A1 => L1_n_106, A2 => y_3(3), B1 => L1_n_70, B2 => L1_n_134, ZN => L1_n_324);
  L1_g29313 : MAOI22D0BWP7T port map(A1 => L1_n_100, A2 => y_0(5), B1 => L1_n_119, B2 => L1_n_61, ZN => L1_n_323);
  L1_g29314 : MAOI22D0BWP7T port map(A1 => L1_n_85, A2 => y_2(0), B1 => L1_n_50, B2 => L1_n_153, ZN => L1_n_322);
  L1_g29315 : MAOI22D0BWP7T port map(A1 => L1_n_100, A2 => y_0(3), B1 => L1_n_136, B2 => L1_n_61, ZN => L1_n_321);
  L1_g29316 : MAOI22D0BWP7T port map(A1 => L1_n_100, A2 => x_0(5), B1 => L1_n_135, B2 => L1_n_47, ZN => L1_n_320);
  L1_g29317 : MAOI22D0BWP7T port map(A1 => L1_n_100, A2 => y_0(0), B1 => L1_n_120, B2 => L1_n_61, ZN => L1_n_319);
  L1_g29318 : MAOI22D0BWP7T port map(A1 => L1_n_100, A2 => y_0(2), B1 => L1_n_142, B2 => L1_n_69, ZN => L1_n_318);
  L1_g29319 : AOI22D0BWP7T port map(A1 => L1_n_85, A2 => x_2(7), B1 => L1_n_99, B2 => x_15(7), ZN => L1_n_317);
  L1_g29320 : OR2D1BWP7T port map(A1 => L1_n_155, A2 => L1_n_59, Z => L1_n_316);
  L1_g29321 : ND4D0BWP7T port map(A1 => L1_n_80, A2 => L1_n_79, A3 => L1_n_78, A4 => L1_n_77, ZN => L1_n_315);
  L1_g29322 : AOI22D0BWP7T port map(A1 => L1_n_103, A2 => y_6(1), B1 => L1_n_90, B2 => y_5(1), ZN => L1_n_314);
  L1_g29323 : AOI22D0BWP7T port map(A1 => L1_n_101, A2 => y_4(1), B1 => L1_n_92, B2 => y_3(1), ZN => L1_n_313);
  L1_g29324 : AOI22D0BWP7T port map(A1 => L1_n_93, A2 => y_9(1), B1 => L1_n_94, B2 => y_13(1), ZN => L1_n_312);
  L1_g29325 : AOI22D0BWP7T port map(A1 => L1_n_82, A2 => y_8(1), B1 => L1_n_83, B2 => y_12(1), ZN => L1_n_311);
  L1_g29326 : AOI22D0BWP7T port map(A1 => L1_n_83, A2 => x_12(1), B1 => L1_n_87, B2 => x_10(1), ZN => L1_n_310);
  L1_g29327 : AOI22D0BWP7T port map(A1 => L1_n_101, A2 => x_4(1), B1 => L1_n_86, B2 => x_14(1), ZN => L1_n_309);
  L1_g29328 : AOI22D0BWP7T port map(A1 => L1_n_93, A2 => y_9(5), B1 => L1_n_94, B2 => y_13(5), ZN => L1_n_308);
  L1_g29329 : AOI22D0BWP7T port map(A1 => L1_n_106, A2 => y_3(1), B1 => L1_n_102, B2 => y_14(1), ZN => L1_n_307);
  L1_g29330 : AOI22D0BWP7T port map(A1 => L1_n_93, A2 => x_9(1), B1 => L1_n_91, B2 => x_7(1), ZN => L1_n_306);
  L1_g29331 : AOI22D0BWP7T port map(A1 => L1_n_88, A2 => x_1(1), B1 => L1_n_90, B2 => x_5(1), ZN => L1_n_305);
  L1_g29332 : AOI22D0BWP7T port map(A1 => L1_n_107, A2 => x_11(8), B1 => L1_n_108, B2 => x_7(8), ZN => L1_n_304);
  L1_g29333 : AOI22D0BWP7T port map(A1 => L1_n_103, A2 => x_6(0), B1 => L1_n_87, B2 => x_10(0), ZN => L1_n_303);
  L1_g29334 : AOI22D0BWP7T port map(A1 => L1_n_81, A2 => x_10(8), B1 => L1_n_99, B2 => x_15(8), ZN => L1_n_302);
  L1_g29335 : AOI22D0BWP7T port map(A1 => L1_n_82, A2 => x_8(0), B1 => L1_n_86, B2 => x_14(0), ZN => L1_n_301);
  L1_g29336 : AOI22D0BWP7T port map(A1 => L1_n_89, A2 => x_9(8), B1 => L1_n_110, B2 => x_13(8), ZN => L1_n_300);
  L1_g29337 : AOI22D0BWP7T port map(A1 => L1_n_92, A2 => x_3(0), B1 => L1_n_91, B2 => x_7(0), ZN => L1_n_299);
  L1_g29338 : AOI22D0BWP7T port map(A1 => L1_n_95, A2 => x_1(8), B1 => L1_n_96, B2 => x_5(8), ZN => L1_n_298);
  L1_g29339 : AOI22D0BWP7T port map(A1 => L1_n_109, A2 => y_8(2), B1 => L1_n_105, B2 => y_12(2), ZN => L1_n_297);
  L1_g29340 : AOI22D0BWP7T port map(A1 => L1_n_88, A2 => x_1(0), B1 => L1_n_90, B2 => x_5(0), ZN => L1_n_296);
  L1_g29341 : AOI22D0BWP7T port map(A1 => L1_n_105, A2 => y_12(8), B1 => L1_n_81, B2 => y_10(8), ZN => L1_n_295);
  L1_g29342 : AOI22D0BWP7T port map(A1 => L1_n_112, A2 => y_4(8), B1 => L1_n_102, B2 => y_14(8), ZN => L1_n_294);
  L1_g29343 : AOI22D0BWP7T port map(A1 => L1_n_83, A2 => x_12(8), B1 => L1_n_87, B2 => x_10(8), ZN => L1_n_293);
  L1_g29344 : AOI22D0BWP7T port map(A1 => L1_n_101, A2 => x_4(8), B1 => L1_n_86, B2 => x_14(8), ZN => L1_n_292);
  L1_g29345 : AOI22D0BWP7T port map(A1 => L1_n_89, A2 => y_9(8), B1 => L1_n_110, B2 => y_13(8), ZN => L1_n_291);
  L1_g29346 : AOI22D0BWP7T port map(A1 => L1_n_106, A2 => y_3(8), B1 => L1_n_108, B2 => y_7(8), ZN => L1_n_290);
  L1_g29347 : AOI22D0BWP7T port map(A1 => L1_n_92, A2 => x_3(8), B1 => L1_n_91, B2 => x_7(8), ZN => L1_n_289);
  L1_g29348 : AOI22D0BWP7T port map(A1 => L1_n_88, A2 => x_1(5), B1 => L1_n_90, B2 => x_5(5), ZN => L1_n_288);
  L1_g29349 : AOI22D0BWP7T port map(A1 => L1_n_106, A2 => x_3(6), B1 => L1_n_89, B2 => x_9(6), ZN => L1_n_287);
  L1_g29350 : AOI22D0BWP7T port map(A1 => L1_n_112, A2 => x_4(6), B1 => L1_n_108, B2 => x_7(6), ZN => L1_n_286);
  L1_g29351 : AOI22D0BWP7T port map(A1 => L1_n_88, A2 => x_1(8), B1 => L1_n_90, B2 => x_5(8), ZN => L1_n_285);
  L1_g29352 : AOI22D0BWP7T port map(A1 => L1_n_107, A2 => x_11(6), B1 => L1_n_99, B2 => x_15(6), ZN => L1_n_284);
  L1_g29353 : AOI22D0BWP7T port map(A1 => L1_n_81, A2 => x_10(6), B1 => L1_n_102, B2 => x_14(6), ZN => L1_n_283);
  L1_g29354 : AOI22D0BWP7T port map(A1 => L1_n_111, A2 => x_0(6), B1 => L1_n_109, B2 => x_8(6), ZN => L1_n_282);
  L1_g29355 : AOI22D0BWP7T port map(A1 => L1_n_82, A2 => y_8(8), B1 => L1_n_103, B2 => y_6(8), ZN => L1_n_281);
  L1_g29356 : AOI22D0BWP7T port map(A1 => L1_n_83, A2 => x_12(4), B1 => L1_n_87, B2 => x_10(4), ZN => L1_n_280);
  L1_g29357 : AOI22D0BWP7T port map(A1 => L1_n_81, A2 => x_10(7), B1 => L1_n_102, B2 => x_14(7), ZN => L1_n_279);
  L1_g29358 : OR2D1BWP7T port map(A1 => L1_n_154, A2 => L1_n_59, Z => L1_n_278);
  L1_g29359 : AOI22D0BWP7T port map(A1 => L1_n_89, A2 => x_9(7), B1 => L1_n_110, B2 => x_13(7), ZN => L1_n_277);
  L1_g29360 : AOI22D0BWP7T port map(A1 => L1_n_82, A2 => x_8(4), B1 => L1_n_103, B2 => x_6(4), ZN => L1_n_276);
  L1_g29361 : AOI22D0BWP7T port map(A1 => L1_n_109, A2 => x_8(7), B1 => L1_n_105, B2 => x_12(7), ZN => L1_n_275);
  L1_g29362 : AOI22D0BWP7T port map(A1 => L1_n_93, A2 => x_9(4), B1 => L1_n_94, B2 => x_13(4), ZN => L1_n_274);
  L1_g29363 : AOI22D0BWP7T port map(A1 => L1_n_88, A2 => x_1(4), B1 => L1_n_90, B2 => x_5(4), ZN => L1_n_273);
  L1_g29364 : AOI22D0BWP7T port map(A1 => L1_n_105, A2 => x_12(5), B1 => L1_n_81, B2 => x_10(5), ZN => L1_n_272);
  L1_g29365 : AOI22D0BWP7T port map(A1 => L1_n_112, A2 => x_4(5), B1 => L1_n_102, B2 => x_14(5), ZN => L1_n_271);
  L1_g29366 : AOI22D0BWP7T port map(A1 => L1_n_89, A2 => x_9(5), B1 => L1_n_110, B2 => x_13(5), ZN => L1_n_270);
  L1_g29367 : AOI22D0BWP7T port map(A1 => L1_n_95, A2 => x_1(5), B1 => L1_n_96, B2 => x_5(5), ZN => L1_n_269);
  L1_g29368 : AOI22D0BWP7T port map(A1 => L1_n_83, A2 => x_12(3), B1 => L1_n_87, B2 => x_10(3), ZN => L1_n_268);
  L1_g29369 : AOI22D0BWP7T port map(A1 => L1_n_81, A2 => x_10(4), B1 => L1_n_102, B2 => x_14(4), ZN => L1_n_267);
  L1_g29370 : AOI22D0BWP7T port map(A1 => L1_n_82, A2 => x_8(3), B1 => L1_n_103, B2 => x_6(3), ZN => L1_n_266);
  L1_g29371 : AOI22D0BWP7T port map(A1 => L1_n_85, A2 => x_2(4), B1 => L1_n_99, B2 => x_15(4), ZN => L1_n_265);
  L1_g29372 : AOI22D0BWP7T port map(A1 => L1_n_93, A2 => x_9(3), B1 => L1_n_91, B2 => x_7(3), ZN => L1_n_264);
  L1_g29373 : AOI22D0BWP7T port map(A1 => L1_n_89, A2 => x_9(4), B1 => L1_n_110, B2 => x_13(4), ZN => L1_n_263);
  L1_g29374 : AOI22D0BWP7T port map(A1 => L1_n_109, A2 => x_8(4), B1 => L1_n_105, B2 => x_12(4), ZN => L1_n_262);
  L1_g29375 : AOI22D0BWP7T port map(A1 => L1_n_88, A2 => x_1(3), B1 => L1_n_90, B2 => x_5(3), ZN => L1_n_261);
  L1_g29376 : AOI22D0BWP7T port map(A1 => L1_n_105, A2 => x_12(3), B1 => L1_n_81, B2 => x_10(3), ZN => L1_n_260);
  L1_g29377 : AOI22D0BWP7T port map(A1 => L1_n_112, A2 => x_4(3), B1 => L1_n_102, B2 => x_14(3), ZN => L1_n_259);
  L1_g29378 : AOI22D0BWP7T port map(A1 => L1_n_83, A2 => x_12(7), B1 => L1_n_87, B2 => x_10(7), ZN => L1_n_258);
  L1_g29379 : AOI22D0BWP7T port map(A1 => L1_n_82, A2 => x_8(7), B1 => L1_n_103, B2 => x_6(7), ZN => L1_n_257);
  L1_g29380 : AOI22D0BWP7T port map(A1 => L1_n_89, A2 => x_9(3), B1 => L1_n_110, B2 => x_13(3), ZN => L1_n_256);
  L1_g29381 : AOI22D0BWP7T port map(A1 => L1_n_95, A2 => x_1(3), B1 => L1_n_96, B2 => x_5(3), ZN => L1_n_255);
  L1_g29382 : AOI22D0BWP7T port map(A1 => L1_n_93, A2 => x_9(7), B1 => L1_n_91, B2 => x_7(7), ZN => L1_n_254);
  L1_g29383 : AOI22D0BWP7T port map(A1 => L1_n_88, A2 => x_1(7), B1 => L1_n_90, B2 => x_5(7), ZN => L1_n_253);
  L1_g29384 : AOI22D0BWP7T port map(A1 => L1_n_102, A2 => x_14(2), B1 => L1_n_108, B2 => x_7(2), ZN => L1_n_252);
  L1_g29385 : AOI22D0BWP7T port map(A1 => L1_n_81, A2 => x_10(2), B1 => L1_n_107, B2 => x_11(2), ZN => L1_n_251);
  L1_g29386 : AOI22D0BWP7T port map(A1 => L1_n_89, A2 => x_9(2), B1 => L1_n_110, B2 => x_13(2), ZN => L1_n_250);
  L1_g29387 : AOI22D0BWP7T port map(A1 => L1_n_109, A2 => x_8(2), B1 => L1_n_105, B2 => x_12(2), ZN => L1_n_249);
  L1_g29388 : AOI22D0BWP7T port map(A1 => L1_n_83, A2 => x_12(6), B1 => L1_n_87, B2 => x_10(6), ZN => L1_n_248);
  L1_g29389 : AOI22D0BWP7T port map(A1 => L1_n_82, A2 => x_8(6), B1 => L1_n_103, B2 => x_6(6), ZN => L1_n_247);
  L1_g29390 : AOI22D0BWP7T port map(A1 => L1_n_81, A2 => x_10(1), B1 => L1_n_102, B2 => x_14(1), ZN => L1_n_246);
  L1_g29391 : AOI22D0BWP7T port map(A1 => L1_n_85, A2 => x_2(1), B1 => L1_n_99, B2 => x_15(1), ZN => L1_n_245);
  L1_g29392 : AOI22D0BWP7T port map(A1 => L1_n_89, A2 => x_9(1), B1 => L1_n_110, B2 => x_13(1), ZN => L1_n_244);
  L1_g29393 : AOI22D0BWP7T port map(A1 => L1_n_95, A2 => x_1(1), B1 => L1_n_96, B2 => x_5(1), ZN => L1_n_243);
  L1_g29394 : AOI22D0BWP7T port map(A1 => L1_n_93, A2 => x_9(6), B1 => L1_n_91, B2 => x_7(6), ZN => L1_n_242);
  L1_g29395 : AOI22D0BWP7T port map(A1 => L1_n_88, A2 => x_1(6), B1 => L1_n_90, B2 => x_5(6), ZN => L1_n_241);
  L1_g29396 : AOI22D0BWP7T port map(A1 => L1_n_109, A2 => x_8(0), B1 => L1_n_81, B2 => x_10(0), ZN => L1_n_240);
  L1_g29397 : AOI22D0BWP7T port map(A1 => L1_n_82, A2 => x_8(2), B1 => L1_n_83, B2 => x_12(2), ZN => L1_n_239);
  L1_g29398 : AOI22D0BWP7T port map(A1 => L1_n_89, A2 => y_9(7), B1 => L1_n_110, B2 => y_13(7), ZN => L1_n_238);
  L1_g29399 : AOI22D0BWP7T port map(A1 => L1_n_89, A2 => x_9(0), B1 => L1_n_110, B2 => x_13(0), ZN => L1_n_237);
  L1_g29400 : AOI22D0BWP7T port map(A1 => L1_n_106, A2 => x_3(0), B1 => L1_n_108, B2 => x_7(0), ZN => L1_n_236);
  L1_g29401 : AOI22D0BWP7T port map(A1 => L1_n_103, A2 => y_6(7), B1 => L1_n_87, B2 => y_10(7), ZN => L1_n_235);
  L1_g29402 : AOI22D0BWP7T port map(A1 => L1_n_82, A2 => y_8(7), B1 => L1_n_86, B2 => y_14(7), ZN => L1_n_234);
  L1_g29403 : AOI22D0BWP7T port map(A1 => L1_n_103, A2 => y_6(5), B1 => L1_n_90, B2 => y_5(5), ZN => L1_n_233);
  L1_g29404 : AOI22D0BWP7T port map(A1 => L1_n_92, A2 => y_3(7), B1 => L1_n_91, B2 => y_7(7), ZN => L1_n_232);
  L1_g29405 : AOI22D0BWP7T port map(A1 => L1_n_111, A2 => y_0(6), B1 => L1_n_102, B2 => y_14(6), ZN => L1_n_231);
  L1_g29406 : AOI22D0BWP7T port map(A1 => L1_n_105, A2 => y_12(6), B1 => L1_n_99, B2 => y_15(6), ZN => L1_n_230);
  L1_g29407 : AOI22D0BWP7T port map(A1 => L1_n_88, A2 => y_1(7), B1 => L1_n_90, B2 => y_5(7), ZN => L1_n_229);
  L1_g29408 : AOI22D0BWP7T port map(A1 => L1_n_89, A2 => y_9(6), B1 => L1_n_110, B2 => y_13(6), ZN => L1_n_228);
  L1_g29409 : AOI22D0BWP7T port map(A1 => L1_n_112, A2 => y_4(6), B1 => L1_n_106, B2 => y_3(6), ZN => L1_n_227);
  L1_g29410 : AOI22D0BWP7T port map(A1 => L1_n_102, A2 => y_14(7), B1 => L1_n_107, B2 => y_11(7), ZN => L1_n_226);
  L1_g29411 : AOI22D0BWP7T port map(A1 => L1_n_106, A2 => y_3(7), B1 => L1_n_99, B2 => y_15(7), ZN => L1_n_225);
  L1_g29412 : AOI22D0BWP7T port map(A1 => L1_n_103, A2 => y_6(6), B1 => L1_n_90, B2 => y_5(6), ZN => L1_n_224);
  L1_g29413 : AOI22D0BWP7T port map(A1 => L1_n_109, A2 => y_8(7), B1 => L1_n_105, B2 => y_12(7), ZN => L1_n_223);
  L1_g29414 : AOI22D0BWP7T port map(A1 => L1_n_88, A2 => y_1(6), B1 => L1_n_91, B2 => y_7(6), ZN => L1_n_222);
  L1_g29415 : AOI22D0BWP7T port map(A1 => L1_n_105, A2 => y_12(5), B1 => L1_n_81, B2 => y_10(5), ZN => L1_n_221);
  L1_g29416 : AOI22D0BWP7T port map(A1 => L1_n_93, A2 => y_9(6), B1 => L1_n_94, B2 => y_13(6), ZN => L1_n_220);
  L1_g29417 : AOI22D0BWP7T port map(A1 => L1_n_82, A2 => y_8(6), B1 => L1_n_83, B2 => y_12(6), ZN => L1_n_219);
  L1_g29418 : AOI22D0BWP7T port map(A1 => L1_n_106, A2 => y_3(5), B1 => L1_n_108, B2 => y_7(5), ZN => L1_n_218);
  L1_g29419 : AOI22D0BWP7T port map(A1 => L1_n_105, A2 => y_12(4), B1 => L1_n_81, B2 => y_10(4), ZN => L1_n_217);
  L1_g29420 : AOI22D0BWP7T port map(A1 => L1_n_109, A2 => y_8(4), B1 => L1_n_112, B2 => y_4(4), ZN => L1_n_216);
  L1_g29421 : AOI22D0BWP7T port map(A1 => L1_n_83, A2 => y_12(8), B1 => L1_n_87, B2 => y_10(8), ZN => L1_n_215);
  L1_g29422 : AOI22D0BWP7T port map(A1 => L1_n_106, A2 => y_3(4), B1 => L1_n_108, B2 => y_7(4), ZN => L1_n_214);
  L1_g29423 : AOI22D0BWP7T port map(A1 => L1_n_95, A2 => y_1(4), B1 => L1_n_96, B2 => y_5(4), ZN => L1_n_213);
  L1_g29424 : AOI22D0BWP7T port map(A1 => L1_n_92, A2 => y_3(8), B1 => L1_n_91, B2 => y_7(8), ZN => L1_n_212);
  L1_g29425 : AOI22D0BWP7T port map(A1 => L1_n_100, A2 => y_0(8), B1 => L1_n_104, B2 => y_2(8), ZN => L1_n_211);
  L1_g29426 : AOI22D0BWP7T port map(A1 => L1_n_102, A2 => y_14(3), B1 => L1_n_108, B2 => y_7(3), ZN => L1_n_210);
  L1_g29427 : AOI22D0BWP7T port map(A1 => L1_n_81, A2 => y_10(3), B1 => L1_n_107, B2 => y_11(3), ZN => L1_n_209);
  L1_g29428 : AOI22D0BWP7T port map(A1 => L1_n_93, A2 => y_9(8), B1 => L1_n_97, B2 => y_11(8), ZN => L1_n_208);
  L1_g29429 : AOI22D0BWP7T port map(A1 => L1_n_89, A2 => y_9(3), B1 => L1_n_110, B2 => y_13(3), ZN => L1_n_207);
  L1_g29430 : AOI22D0BWP7T port map(A1 => L1_n_95, A2 => y_1(3), B1 => L1_n_96, B2 => y_5(3), ZN => L1_n_206);
  L1_g29431 : AOI22D0BWP7T port map(A1 => L1_n_112, A2 => y_4(5), B1 => L1_n_102, B2 => y_14(5), ZN => L1_n_205);
  L1_g29432 : AOI22D0BWP7T port map(A1 => L1_n_89, A2 => y_9(5), B1 => L1_n_110, B2 => y_13(5), ZN => L1_n_204);
  L1_g29433 : AOI22D0BWP7T port map(A1 => L1_n_106, A2 => y_3(2), B1 => L1_n_102, B2 => y_14(2), ZN => L1_n_203);
  L1_g29434 : AOI22D0BWP7T port map(A1 => L1_n_81, A2 => y_10(2), B1 => L1_n_84, B2 => y_6(2), ZN => L1_n_202);
  L1_g29435 : AOI22D0BWP7T port map(A1 => L1_n_88, A2 => y_1(5), B1 => L1_n_91, B2 => y_7(5), ZN => L1_n_201);
  L1_g29436 : AOI22D0BWP7T port map(A1 => L1_n_89, A2 => y_9(2), B1 => L1_n_110, B2 => y_13(2), ZN => L1_n_200);
  L1_g29437 : AOI22D0BWP7T port map(A1 => L1_n_95, A2 => y_1(2), B1 => L1_n_96, B2 => y_5(2), ZN => L1_n_199);
  L1_g29438 : AOI22D0BWP7T port map(A1 => L1_n_111, A2 => y_0(2), B1 => L1_n_112, B2 => y_4(2), ZN => L1_n_198);
  L1_g29439 : AOI22D0BWP7T port map(A1 => L1_n_82, A2 => y_8(5), B1 => L1_n_83, B2 => y_12(5), ZN => L1_n_197);
  L1_g29440 : AOI22D0BWP7T port map(A1 => L1_n_81, A2 => y_10(1), B1 => L1_n_84, B2 => y_6(1), ZN => L1_n_196);
  L1_g29441 : AOI22D0BWP7T port map(A1 => L1_n_107, A2 => y_11(1), B1 => L1_n_108, B2 => y_7(1), ZN => L1_n_195);
  L1_g29442 : AOI22D0BWP7T port map(A1 => L1_n_89, A2 => y_9(1), B1 => L1_n_110, B2 => y_13(1), ZN => L1_n_194);
  L1_g29443 : AOI22D0BWP7T port map(A1 => L1_n_109, A2 => y_8(1), B1 => L1_n_105, B2 => y_12(1), ZN => L1_n_193);
  L1_g29444 : AOI22D0BWP7T port map(A1 => L1_n_111, A2 => y_0(1), B1 => L1_n_112, B2 => y_4(1), ZN => L1_n_192);
  L1_g29445 : AOI22D0BWP7T port map(A1 => L1_n_94, A2 => x_13(5), B1 => L1_n_97, B2 => x_11(5), ZN => L1_n_191);
  L1_g29446 : AOI22D0BWP7T port map(A1 => L1_n_103, A2 => y_6(4), B1 => L1_n_87, B2 => y_10(4), ZN => L1_n_190);
  L1_g29447 : AOI22D0BWP7T port map(A1 => L1_n_107, A2 => y_11(0), B1 => L1_n_108, B2 => y_7(0), ZN => L1_n_189);
  L1_g29448 : AOI22D0BWP7T port map(A1 => L1_n_81, A2 => y_10(0), B1 => L1_n_99, B2 => y_15(0), ZN => L1_n_188);
  L1_g29449 : AOI22D0BWP7T port map(A1 => L1_n_82, A2 => y_8(4), B1 => L1_n_86, B2 => y_14(4), ZN => L1_n_187);
  L1_g29450 : AOI22D0BWP7T port map(A1 => L1_n_95, A2 => y_1(0), B1 => L1_n_96, B2 => y_5(0), ZN => L1_n_186);
  L1_g29451 : AOI22D0BWP7T port map(A1 => L1_n_109, A2 => y_8(0), B1 => L1_n_105, B2 => y_12(0), ZN => L1_n_185);
  L1_g29452 : AOI22D0BWP7T port map(A1 => L1_n_103, A2 => x_6(5), B1 => L1_n_93, B2 => x_9(5), ZN => L1_n_184);
  L1_g29453 : AOI22D0BWP7T port map(A1 => L1_n_100, A2 => y_0(4), B1 => L1_n_104, B2 => y_2(4), ZN => L1_n_183);
  L1_g29454 : AOI22D0BWP7T port map(A1 => L1_n_92, A2 => y_3(4), B1 => L1_n_91, B2 => y_7(4), ZN => L1_n_182);
  L1_g29455 : AOI22D0BWP7T port map(A1 => L1_n_95, A2 => y_1(1), B1 => L1_n_96, B2 => y_5(1), ZN => L1_n_181);
  L1_g29456 : AOI22D0BWP7T port map(A1 => L1_n_93, A2 => y_9(4), B1 => L1_n_97, B2 => y_11(4), ZN => L1_n_180);
  L1_g29457 : AOI22D0BWP7T port map(A1 => L1_n_101, A2 => y_4(0), B1 => L1_n_91, B2 => y_7(0), ZN => L1_n_179);
  L1_g29458 : AOI22D0BWP7T port map(A1 => L1_n_103, A2 => y_6(3), B1 => L1_n_87, B2 => y_10(3), ZN => L1_n_178);
  L1_g29459 : AOI22D0BWP7T port map(A1 => L1_n_82, A2 => y_8(3), B1 => L1_n_86, B2 => y_14(3), ZN => L1_n_177);
  L1_g29460 : AOI22D0BWP7T port map(A1 => L1_n_82, A2 => x_8(5), B1 => L1_n_83, B2 => x_12(5), ZN => L1_n_176);
  L1_g29461 : AOI22D0BWP7T port map(A1 => L1_n_90, A2 => y_5(0), B1 => L1_n_92, B2 => y_3(0), ZN => L1_n_175);
  L1_g29462 : AOI22D0BWP7T port map(A1 => L1_n_93, A2 => y_9(3), B1 => L1_n_91, B2 => y_7(3), ZN => L1_n_174);
  L1_g29463 : AOI22D0BWP7T port map(A1 => L1_n_88, A2 => y_1(3), B1 => L1_n_90, B2 => y_5(3), ZN => L1_n_173);
  L1_g29464 : AOI22D0BWP7T port map(A1 => L1_n_107, A2 => y_11(2), B1 => L1_n_108, B2 => y_7(2), ZN => L1_n_172);
  L1_g29465 : AOI22D0BWP7T port map(A1 => L1_n_97, A2 => y_11(0), B1 => L1_n_113, B2 => y_15(0), ZN => L1_n_171);
  L1_g29466 : AOI22D0BWP7T port map(A1 => L1_n_82, A2 => y_8(0), B1 => L1_n_83, B2 => y_12(0), ZN => L1_n_170);
  L1_g29467 : AOI22D0BWP7T port map(A1 => L1_n_93, A2 => x_9(2), B1 => L1_n_113, B2 => x_15(2), ZN => L1_n_169);
  L1_g29468 : AOI22D0BWP7T port map(A1 => L1_n_103, A2 => y_6(2), B1 => L1_n_93, B2 => y_9(2), ZN => L1_n_168);
  L1_g29469 : AOI22D0BWP7T port map(A1 => L1_n_94, A2 => y_13(2), B1 => L1_n_97, B2 => y_11(2), ZN => L1_n_167);
  L1_g29470 : AOI22D0BWP7T port map(A1 => L1_n_109, A2 => y_8(6), B1 => L1_n_107, B2 => y_11(6), ZN => L1_n_166);
  L1_g29471 : AOI22D0BWP7T port map(A1 => L1_n_103, A2 => x_6(2), B1 => L1_n_97, B2 => x_11(2), ZN => L1_n_165);
  L1_g29472 : AOI22D0BWP7T port map(A1 => L1_n_92, A2 => y_3(2), B1 => L1_n_91, B2 => y_7(2), ZN => L1_n_164);
  L1_g29473 : AOI22D0BWP7T port map(A1 => L1_n_88, A2 => y_1(2), B1 => L1_n_90, B2 => y_5(2), ZN => L1_n_163);
  L1_g29474 : AOI22D0BWP7T port map(A1 => L1_n_88, A2 => x_1(2), B1 => L1_n_90, B2 => x_5(2), ZN => L1_n_162);
  L1_g29475 : AOI22D0BWP7T port map(A1 => L1_n_111, A2 => x_0(0), B1 => L1_n_102, B2 => x_14(0), ZN => L1_n_161);
  L1_g29476 : INVD1BWP7T port map(I => L1_n_156, ZN => L1_n_157);
  L1_g29477 : AOI22D0BWP7T port map(A1 => L1_n_55, A2 => y_9(0), B1 => L1_n_53, B2 => y_13(0), ZN => L1_n_153);
  L1_g29478 : CKND2D0BWP7T port map(A1 => L1_n_85, A2 => y_2(6), ZN => L1_n_152);
  L1_g29479 : AO22D0BWP7T port map(A1 => L1_n_51, A2 => y_1(4), B1 => y_5(4), B2 => L1_n_66, Z => L1_n_151);
  L1_g29480 : CKND2D0BWP7T port map(A1 => L1_n_95, A2 => x_1(6), ZN => L1_n_150);
  L1_g29481 : AOI22D0BWP7T port map(A1 => L1_n_55, A2 => y_9(4), B1 => L1_n_53, B2 => y_13(4), ZN => L1_n_149);
  L1_g29482 : AOI22D0BWP7T port map(A1 => L1_n_51, A2 => y_9(7), B1 => L1_n_66, B2 => y_13(7), ZN => L1_n_148);
  L1_g29483 : AO22D0BWP7T port map(A1 => L1_n_51, A2 => y_1(8), B1 => y_5(8), B2 => L1_n_66, Z => L1_n_147);
  L1_g29484 : AOI22D0BWP7T port map(A1 => L1_n_43, A2 => y_11(1), B1 => L1_n_63, B2 => y_15(1), ZN => L1_n_146);
  L1_g29485 : OAI21D0BWP7T port map(A1 => L1_n_57, A2 => count_1_s(1), B => enable_s, ZN => L1_n_145);
  L1_g29486 : AOI22D0BWP7T port map(A1 => L1_n_43, A2 => x_11(7), B1 => L1_n_63, B2 => x_15(7), ZN => L1_n_144);
  L1_g29487 : AOI22D0BWP7T port map(A1 => L1_n_43, A2 => x_3(2), B1 => L1_n_63, B2 => x_7(2), ZN => L1_n_143);
  L1_g29488 : AOI22D0BWP7T port map(A1 => L1_n_43, A2 => y_10(2), B1 => L1_n_63, B2 => y_14(2), ZN => L1_n_142);
  L1_g29489 : AOI22D0BWP7T port map(A1 => L1_n_45, A2 => x_1(4), B1 => L1_n_49, B2 => x_5(4), ZN => L1_n_141);
  L1_g29490 : ND2D1BWP7T port map(A1 => L1_n_118, A2 => L1_n_73, ZN => L1_n_160);
  L1_g29491 : ND3D0BWP7T port map(A1 => L1_n_72, A2 => L1_n_76, A3 => L1_n_18, ZN => L1_n_159);
  L1_g29492 : NR3D0BWP7T port map(A1 => L1_n_73, A2 => L1_n_75, A3 => L1_state(0), ZN => L1_n_158);
  L1_g29493 : NR3D0BWP7T port map(A1 => L1_n_73, A2 => L1_n_74, A3 => L1_state(0), ZN => L1_n_156);
  L1_g29496 : IND2D1BWP7T port map(A1 => L1_n_72, B1 => L1_n_118, ZN => L1_n_155);
  L1_g29497 : OR2D1BWP7T port map(A1 => L1_n_117, A2 => L1_n_72, Z => L1_n_154);
  L1_g29498 : AOI22D0BWP7T port map(A1 => L1_n_45, A2 => x_3(3), B1 => L1_n_49, B2 => x_7(3), ZN => L1_n_140);
  L1_g29499 : AOI22D0BWP7T port map(A1 => L1_n_51, A2 => x_9(0), B1 => L1_n_66, B2 => x_13(0), ZN => L1_n_139);
  L1_g29500 : AOI22D0BWP7T port map(A1 => L1_n_43, A2 => x_11(3), B1 => L1_n_63, B2 => x_15(3), ZN => L1_n_138);
  L1_g29501 : AOI22D0BWP7T port map(A1 => L1_n_45, A2 => y_1(8), B1 => L1_n_49, B2 => y_5(8), ZN => L1_n_137);
  L1_g29502 : AOI22D0BWP7T port map(A1 => L1_n_43, A2 => y_11(3), B1 => L1_n_63, B2 => y_15(3), ZN => L1_n_136);
  L1_g29503 : AOI22D0BWP7T port map(A1 => L1_n_43, A2 => x_3(5), B1 => L1_n_63, B2 => x_7(5), ZN => L1_n_135);
  L1_g29504 : AOI22D0BWP7T port map(A1 => L1_n_55, A2 => y_8(3), B1 => L1_n_53, B2 => y_12(3), ZN => L1_n_134);
  L1_g29505 : AOI22D0BWP7T port map(A1 => L1_n_45, A2 => x_1(7), B1 => L1_n_49, B2 => x_5(7), ZN => L1_n_133);
  L1_g29506 : AOI22D0BWP7T port map(A1 => L1_n_43, A2 => x_3(4), B1 => L1_n_63, B2 => x_7(4), ZN => L1_n_132);
  L1_g29507 : AOI22D0BWP7T port map(A1 => L1_n_45, A2 => x_1(2), B1 => L1_n_49, B2 => x_5(2), ZN => L1_n_131);
  L1_g29508 : AOI22D0BWP7T port map(A1 => L1_n_43, A2 => x_11(6), B1 => L1_n_63, B2 => x_15(6), ZN => L1_n_130);
  L1_g29509 : AOI22D0BWP7T port map(A1 => L1_n_45, A2 => x_0(8), B1 => L1_n_49, B2 => x_4(8), ZN => L1_n_129);
  L1_g29510 : AOI22D0BWP7T port map(A1 => L1_n_45, A2 => y_1(7), B1 => L1_n_49, B2 => y_5(7), ZN => L1_n_128);
  L1_g29511 : AOI22D0BWP7T port map(A1 => L1_n_55, A2 => x_11(5), B1 => L1_n_53, B2 => x_15(5), ZN => L1_n_127);
  L1_g29512 : AOI22D0BWP7T port map(A1 => L1_n_45, A2 => x_1(0), B1 => L1_n_49, B2 => x_5(0), ZN => L1_n_126);
  L1_g29513 : AOI22D0BWP7T port map(A1 => L1_n_43, A2 => x_11(1), B1 => L1_n_63, B2 => x_15(1), ZN => L1_n_125);
  L1_g29514 : AOI22D0BWP7T port map(A1 => L1_n_51, A2 => x_9(8), B1 => L1_n_66, B2 => x_13(8), ZN => L1_n_124);
  L1_g29515 : AOI22D0BWP7T port map(A1 => L1_n_45, A2 => x_0(1), B1 => L1_n_49, B2 => x_4(1), ZN => L1_n_123);
  L1_g29516 : AOI22D0BWP7T port map(A1 => L1_n_43, A2 => y_11(6), B1 => L1_n_63, B2 => y_15(6), ZN => L1_n_122);
  L1_g29517 : AOI22D0BWP7T port map(A1 => L1_n_45, A2 => y_1(5), B1 => L1_n_49, B2 => y_5(5), ZN => L1_n_121);
  L1_g29518 : AOI22D0BWP7T port map(A1 => L1_n_51, A2 => y_9(0), B1 => L1_n_66, B2 => y_13(0), ZN => L1_n_120);
  L1_g29519 : AOI22D0BWP7T port map(A1 => L1_n_43, A2 => y_11(5), B1 => L1_n_63, B2 => y_15(5), ZN => L1_n_119);
  L1_g29521 : INVD0BWP7T port map(I => L1_n_99, ZN => L1_n_98);
  L1_g29522 : ND2D1BWP7T port map(A1 => L1_n_74, A2 => L1_n_35, ZN => L1_n_118);
  L1_g29523 : NR2D1BWP7T port map(A1 => L1_n_76, A2 => FE_OFN0_reset, ZN => L1_n_117);
  L1_g29524 : NR2XD0BWP7T port map(A1 => L1_n_68, A2 => FE_OFN0_reset, ZN => L1_n_116);
  L1_g29525 : NR2XD0BWP7T port map(A1 => L1_n_60, A2 => FE_OFN0_reset, ZN => L1_n_115);
  L1_g29526 : NR2XD0BWP7T port map(A1 => L1_n_46, A2 => FE_OFN0_reset, ZN => L1_n_114);
  L1_g29527 : NR2D1BWP7T port map(A1 => L1_n_61, A2 => L1_n_62, ZN => L1_n_113);
  L1_g29528 : NR2D1P5BWP7T port map(A1 => L1_n_48, A2 => L1_n_70, ZN => L1_n_112);
  L1_g29529 : NR2D1P5BWP7T port map(A1 => L1_n_44, A2 => L1_n_70, ZN => L1_n_111);
  L1_g29530 : NR2D1P5BWP7T port map(A1 => L1_n_50, A2 => L1_n_54, ZN => L1_n_110);
  L1_g29531 : INR2D2BWP7T port map(A1 => L1_n_55, B1 => L1_n_70, ZN => L1_n_109);
  L1_g29532 : NR2D1P5BWP7T port map(A1 => L1_n_48, A2 => L1_n_56, ZN => L1_n_108);
  L1_g29533 : INR2D2BWP7T port map(A1 => L1_n_55, B1 => L1_n_56, ZN => L1_n_107);
  L1_g29534 : NR2D1P5BWP7T port map(A1 => L1_n_44, A2 => L1_n_56, ZN => L1_n_106);
  L1_g29535 : NR2D1P5BWP7T port map(A1 => L1_n_70, A2 => L1_n_54, ZN => L1_n_105);
  L1_g29536 : NR2D1P5BWP7T port map(A1 => L1_n_42, A2 => L1_n_57, ZN => L1_n_104);
  L1_g29537 : NR2D1P5BWP7T port map(A1 => L1_n_62, A2 => L1_n_57, ZN => L1_n_103);
  L1_g29538 : NR2D1P5BWP7T port map(A1 => L1_n_58, A2 => L1_n_54, ZN => L1_n_102);
  L1_g29539 : NR2D1P5BWP7T port map(A1 => L1_n_57, A2 => L1_n_67, ZN => L1_n_101);
  L1_g29540 : NR2D1P5BWP7T port map(A1 => L1_n_52, A2 => L1_n_57, ZN => L1_n_100);
  L1_g29541 : NR2D1P5BWP7T port map(A1 => L1_n_56, A2 => L1_n_54, ZN => L1_n_99);
  L1_g29542 : AOI22D0BWP7T port map(A1 => L1_n_37, A2 => count_1_s(1), B1 => count_2_s(1), B2 => L1_n_36, ZN => L1_n_80);
  L1_g29543 : AOI22D0BWP7T port map(A1 => L1_n_40, A2 => count_1_s(2), B1 => count_2_s(2), B2 => L1_n_39, ZN => L1_n_79);
  L1_g29544 : XNR2D1BWP7T port map(A1 => count_2_s(3), A2 => count_1_s(3), ZN => L1_n_78);
  L1_g29545 : XNR2D1BWP7T port map(A1 => count_2_s(0), A2 => count_1_s(0), ZN => L1_n_77);
  L1_g29546 : NR2D1BWP7T port map(A1 => L1_n_42, A2 => L1_n_61, ZN => L1_n_97);
  L1_g29547 : NR2D1BWP7T port map(A1 => L1_n_48, A2 => L1_n_50, ZN => L1_n_96);
  L1_g29548 : NR2D1BWP7T port map(A1 => L1_n_44, A2 => L1_n_50, ZN => L1_n_95);
  L1_g29549 : NR2D1P5BWP7T port map(A1 => L1_n_61, A2 => L1_n_67, ZN => L1_n_94);
  L1_g29550 : NR2D1BWP7T port map(A1 => L1_n_52, A2 => L1_n_61, ZN => L1_n_93);
  L1_g29551 : NR2D1P5BWP7T port map(A1 => L1_n_42, A2 => L1_n_47, ZN => L1_n_92);
  L1_g29552 : NR2D1P5BWP7T port map(A1 => L1_n_47, A2 => L1_n_62, ZN => L1_n_91);
  L1_g29553 : NR2D1P5BWP7T port map(A1 => L1_n_47, A2 => L1_n_67, ZN => L1_n_90);
  L1_g29554 : INR2D2BWP7T port map(A1 => L1_n_55, B1 => L1_n_50, ZN => L1_n_89);
  L1_g29555 : NR2D1P5BWP7T port map(A1 => L1_n_47, A2 => L1_n_52, ZN => L1_n_88);
  L1_g29556 : NR2D1P5BWP7T port map(A1 => L1_n_42, A2 => L1_n_69, ZN => L1_n_87);
  L1_g29557 : NR2D1P5BWP7T port map(A1 => L1_n_69, A2 => L1_n_62, ZN => L1_n_86);
  L1_g29558 : NR2D1P5BWP7T port map(A1 => L1_n_44, A2 => L1_n_58, ZN => L1_n_85);
  L1_g29559 : NR2D1P5BWP7T port map(A1 => L1_n_48, A2 => L1_n_58, ZN => L1_n_84);
  L1_g29560 : NR2D1P5BWP7T port map(A1 => L1_n_69, A2 => L1_n_67, ZN => L1_n_83);
  L1_g29561 : NR2D1P5BWP7T port map(A1 => L1_n_69, A2 => L1_n_52, ZN => L1_n_82);
  L1_g29562 : INR2D2BWP7T port map(A1 => L1_n_55, B1 => L1_n_58, ZN => L1_n_81);
  L1_g29563 : CKND1BWP7T port map(I => L1_n_75, ZN => L1_n_76);
  L1_g29565 : INVD1BWP7T port map(I => L1_n_69, ZN => L1_n_68);
  L1_g29566 : INVD1BWP7T port map(I => L1_n_67, ZN => L1_n_66);
  L1_g29567 : INVD1BWP7T port map(I => L1_n_65, ZN => L1_n_64);
  L1_g29568 : INVD1BWP7T port map(I => L1_n_63, ZN => L1_n_62);
  L1_g29569 : INVD1BWP7T port map(I => L1_n_61, ZN => L1_n_60);
  L1_g29570 : ND2D1BWP7T port map(A1 => L1_n_39, A2 => enable_s, ZN => L1_n_75);
  L1_g29571 : ND2D1BWP7T port map(A1 => enable_s, A2 => count_1_s(2), ZN => L1_n_74);
  L1_g29572 : ND2D1BWP7T port map(A1 => count_1_s(1), A2 => L1_n_35, ZN => L1_n_73);
  L1_g29573 : NR2XD0BWP7T port map(A1 => count_1_s(1), A2 => FE_OFN0_reset, ZN => L1_n_72);
  L1_g29574 : NR2XD0BWP7T port map(A1 => L1_range_state_out(0), A2 => L1_range_state_out(1), ZN => L1_n_71);
  L1_g29575 : IND2D1BWP7T port map(A1 => count_2_s(0), B1 => L1_n_37, ZN => L1_n_70);
  L1_g29576 : IND2D1BWP7T port map(A1 => count_1_s(0), B1 => count_1_s(3), ZN => L1_n_69);
  L1_g29577 : CKND2D1BWP7T port map(A1 => L1_n_36, A2 => count_1_s(2), ZN => L1_n_67);
  L1_g29578 : ND2D1BWP7T port map(A1 => L1_range_state_out(1), A2 => L1_range_state_out(0), ZN => L1_n_65);
  L1_g29579 : NR2D1BWP7T port map(A1 => L1_n_36, A2 => L1_n_39, ZN => L1_n_63);
  L1_g29580 : CKND2D1BWP7T port map(A1 => count_1_s(3), A2 => count_1_s(0), ZN => L1_n_61);
  L1_g29581 : INVD1BWP7T port map(I => L1_n_54, ZN => L1_n_53);
  L1_g29582 : INVD1BWP7T port map(I => L1_n_52, ZN => L1_n_51);
  L1_g29583 : INVD1BWP7T port map(I => L1_n_49, ZN => L1_n_48);
  L1_g29584 : INVD1BWP7T port map(I => L1_n_47, ZN => L1_n_46);
  L1_g29585 : INVD1BWP7T port map(I => L1_n_45, ZN => L1_n_44);
  L1_g29586 : INVD1BWP7T port map(I => L1_n_43, ZN => L1_n_42);
  L1_g29587 : NR2XD0BWP7T port map(A1 => L1_n_41, A2 => FE_OFN0_reset, ZN => L1_n_59);
  L1_g29588 : IND2D1BWP7T port map(A1 => count_2_s(0), B1 => count_2_s(1), ZN => L1_n_58);
  L1_g29589 : OR2D1BWP7T port map(A1 => count_1_s(0), A2 => count_1_s(3), Z => L1_n_57);
  L1_g29590 : CKND2D1BWP7T port map(A1 => count_2_s(1), A2 => count_2_s(0), ZN => L1_n_56);
  L1_g29591 : INR2D1BWP7T port map(A1 => count_2_s(3), B1 => count_2_s(2), ZN => L1_n_55);
  L1_g29592 : CKND2D1BWP7T port map(A1 => count_2_s(3), A2 => count_2_s(2), ZN => L1_n_54);
  L1_g29593 : CKND2D1BWP7T port map(A1 => L1_n_39, A2 => L1_n_36, ZN => L1_n_52);
  L1_g29594 : ND2D1BWP7T port map(A1 => L1_n_37, A2 => count_2_s(0), ZN => L1_n_50);
  L1_g29595 : NR2D1BWP7T port map(A1 => L1_n_40, A2 => count_2_s(3), ZN => L1_n_49);
  L1_g29596 : IND2D1BWP7T port map(A1 => count_1_s(3), B1 => count_1_s(0), ZN => L1_n_47);
  L1_g29597 : NR2D1BWP7T port map(A1 => count_2_s(2), A2 => count_2_s(3), ZN => L1_n_45);
  L1_g29598 : NR2D1BWP7T port map(A1 => L1_n_36, A2 => count_1_s(2), ZN => L1_n_43);
  L1_g29599 : INVD0BWP7T port map(I => L1_n_702, ZN => L1_n_41);
  L1_g29600 : CKND1BWP7T port map(I => count_2_s(2), ZN => L1_n_40);
  L1_g29601 : INVD1BWP7T port map(I => count_1_s(2), ZN => L1_n_39);
  L1_g29607 : INVD1BWP7T port map(I => count_2_s(1), ZN => L1_n_37);
  L1_g29614 : INVD1BWP7T port map(I => count_1_s(1), ZN => L1_n_36);
  L1_g29615 : INVD0BWP7T port map(I => FE_OFN0_reset, ZN => L1_n_35);
  L1_col_reg_0 : DFD0BWP7T port map(CP => CTS_6, D => L1_n_400, Q => L1_n_19, QN => L1_n_3);
  L1_col_reg_1 : DFD0BWP7T port map(CP => CTS_6, D => L1_n_399, Q => L1_n_20, QN => L1_n_15);
  L1_col_reg_2 : DFD0BWP7T port map(CP => CTS_6, D => L1_n_398, Q => L1_n_21, QN => L1_n_16);
  L1_col_reg_3 : DFD0BWP7T port map(CP => CTS_6, D => L1_n_413, Q => L1_n_22, QN => L1_n_13);
  L1_col_reg_4 : DFD0BWP7T port map(CP => CTS_6, D => L1_n_401, Q => L1_n_23, QN => L1_n_12);
  L1_col_reg_5 : DFD0BWP7T port map(CP => CTS_6, D => L1_n_412, Q => L1_n_24, QN => L1_n_11);
  L1_col_reg_6 : DFD0BWP7T port map(CP => CTS_6, D => L1_n_411, Q => L1_n_25, QN => L1_n_17);
  L1_col_reg_7 : DFD0BWP7T port map(CP => CTS_6, D => L1_n_410, Q => L1_n_26, QN => L1_n_9);
  L1_col_reg_8 : DFD0BWP7T port map(CP => CTS_6, D => L1_n_397, Q => L1_n_27, QN => L1_n_8);
  L1_col_reg_9 : DFD0BWP7T port map(CP => CTS_6, D => L1_n_396, Q => L1_n_28, QN => L1_n_14);
  L1_col_reg_10 : DFD0BWP7T port map(CP => CTS_6, D => L1_n_409, Q => L1_n_29, QN => L1_n_6);
  L1_col_reg_11 : DFD0BWP7T port map(CP => CTS_6, D => L1_n_403, Q => L1_n_30, QN => L1_n_10);
  L1_col_reg_12 : DFD0BWP7T port map(CP => CTS_6, D => L1_n_408, Q => L1_n_31, QN => L1_n_4);
  L1_col_reg_13 : DFD0BWP7T port map(CP => CTS_6, D => L1_n_402, Q => L1_n_32, QN => L1_n_7);
  L1_col_reg_14 : DFD0BWP7T port map(CP => CTS_6, D => L1_n_407, Q => FE_PHN15_L1_n_33, QN => L1_n_5);
  L1_col_reg_15 : DFD0BWP7T port map(CP => CTS_6, D => L1_n_406, Q => L1_n_34, QN => L1_n_2);
  L1_drc_bufs29616 : INVD5BWP7T port map(I => L1_n_17, ZN => col(6));
  L1_drc_bufs29620 : INVD5BWP7T port map(I => L1_n_16, ZN => col(2));
  L1_drc_bufs29624 : INVD5BWP7T port map(I => L1_n_15, ZN => col(1));
  L1_drc_bufs29628 : INVD5BWP7T port map(I => L1_n_14, ZN => col(9));
  L1_drc_bufs29632 : INVD5BWP7T port map(I => L1_n_13, ZN => col(3));
  L1_drc_bufs29636 : INVD5BWP7T port map(I => L1_n_12, ZN => col(4));
  L1_drc_bufs29640 : INVD5BWP7T port map(I => L1_n_11, ZN => col(5));
  L1_drc_bufs29644 : INVD5BWP7T port map(I => L1_n_10, ZN => col(11));
  L1_drc_bufs29648 : INVD5BWP7T port map(I => L1_n_9, ZN => col(7));
  L1_drc_bufs29652 : INVD5BWP7T port map(I => L1_n_8, ZN => col(8));
  L1_drc_bufs29656 : INVD5BWP7T port map(I => L1_n_7, ZN => col(13));
  L1_drc_bufs29660 : INVD5BWP7T port map(I => L1_n_6, ZN => col(10));
  L1_drc_bufs29664 : INVD5BWP7T port map(I => L1_n_5, ZN => col(14));
  L1_drc_bufs29668 : INVD5BWP7T port map(I => L1_n_4, ZN => col(12));
  L1_drc_bufs29672 : INVD5BWP7T port map(I => L1_n_3, ZN => col(0));
  L1_drc_bufs29676 : INVD5BWP7T port map(I => L1_n_2, ZN => col(15));
  L1_g2 : IND2D1BWP7T port map(A1 => L1_n_117, B1 => L1_n_73, ZN => L1_n_1);
  L1_g29711 : INR3D0BWP7T port map(A1 => L1_n_72, B1 => L1_n_74, B2 => L1_state(0), ZN => L1_n_0);
  L1_g29712 : NR3D0BWP7T port map(A1 => L1_n_532, A2 => L1_n_724, A3 => L1_n_71, ZN => L1_n_719);
  L1_g29716 : CKXOR2D1BWP7T port map(A1 => L1_n_552, A2 => L1_n_508, Z => L1_n_723);
  L1_range_state_out_reg_0 : DFKCND1BWP7T port map(CN => L1_n_35, CP => CTS_6, D => L1_n_701, Q => L1_range_state_out(0), QN => L1_n_38);
  L1_g29719 : AOI21D0BWP7T port map(A1 => L1_n_64, A2 => L1_n_569, B => L1_n_553, ZN => L1_n_724);
  L1_g29720 : IAO21D0BWP7T port map(A1 => L1_n_725, A2 => L1_n_554, B => L1_n_517, ZN => L1_n_726);
  L1_g3 : INR2D1BWP7T port map(A1 => L1_n_64, B1 => L1_n_559, ZN => L1_n_725);

end routed;
