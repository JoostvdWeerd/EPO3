library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.numeric_std.ALL;

architecture behaviour of enemy is

signal R1,R2,R3,R4,R5,R6,R7,R8,R9,R10,R11,R12,R13,R14,R15,R16,R17,R18,R19,R20,R21,R22,R23,R24,R25,R26 : std_logic_vector(31 downto 0);
signal G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,G21,G22,G23,G24,G25,G26 : std_logic_vector(31 downto 0);
signal B1,B2,B3,B4,B5,B6,B7,B8,B9,B10,B11,B12,B13,B14,B15,B16,B17,B18,B19,B20,B21,B22,B23,B24,B25,B26 : std_logic_vector(31 downto 0);

begin

-- red sprite definition
R1 <= "00000000000000011111110000000000";
R2 <= "00000000000000011000111100000000";
R3 <= "00000000000001111100001111000000";
R4 <= "00000000000110111111100111100000";
R5 <= "00000000011100110011110001110000";
R6 <= "00000000000001111100011100011000";
R7 <= "00000000011111001111000111001100";
R8 <= "00000000000111100011110001100110";
R9 <= "00000000000001110000111100111010";
R10 <="00000011000001111111001110001111";
R11 <="00000111110001100000000111111111";
R12 <="00001111110000111000111000111111";
R13 <="00011111111100011111000111111110";
R14<= "00011111111100011111000111111110";
R15<= "00001111110000111000111000111111";
R16<= "00000111110001100000000111111111";
R17<= "00000011000001111111001110001111";
R18<= "00000000000001110000111100111010";
R19<= "00000000000111100011110001100110";
R20<= "00000000011111001111000111001100";
R21<= "00000000000001111100011100011000";
R22<= "00000000011100110011110001110000";
R23<= "00000000000110111111100111100000";
R24<= "00000000000001111100001111000000";
R25<= "00000000000000011000111100000000";
R26<= "00000000000000011111110000000000";

-- green sprite definition
G1 <= "00000000000000100000000000000000";
G2 <= "00000000000111100000000000000000";
G3 <= "00000000111110000000000000000000";
G4 <= "00000011111000000000000000000000";
G5 <= "00001111100000000000000000000000";
G6 <= "00111110000000000000000000000000";
G7 <= "01111000000000000000000000000000";
G8 <= "01111111111000000000000000000000";
G9 <= "00000000000000000000000000000000";
G10<= "00000000000000000000000000000000";
G11<= "00000000000000011111111000000000";
G12<= "00000011110000000111000000000000";
G13<= "00000111111111100000000000000000";
G14<= "00000111111111100000000000000000";
G15<= "00000011110000000111000000000000";
G16<= "00000000000000011111111000000000";
G17<= "00000000000000000000000000000000";
G18<= "00000000000000000000000000000000";
G19<= "01111111111000000000000000000000";
G20<= "01111000000000000000000000000000";
G21<= "00111110000000000000000000000000";
G22<= "00001111100000000000000000000000";
G23<= "00000011111000000000000000000000";
G24<= "00000000111110000000000000000000";
G25<= "00000000000111100000000000000000";
G26<= "00000000000000100000000000000000";

-- blue sprite definition
B1 <= "00000000000000000000000000000000";  
B2 <= "00000000000000000000000000000000";
B3 <= "00000000000000000000000000000000";
B4 <= "00000000000000000000000000000000";
B5 <= "00000000000000000000000000000000";
B6 <= "00000000000000000000000000000000";
B7 <= "00000000000000000000000000000000";
B8 <= "00000000000000000000000000000000";
B9 <= "00000000000000000000000000000000";
B10<= "00000000000000000000000000000000";
B11<= "00000000000000000000000000000000";
B12<= "00000000000000000000000000000111";
B13<= "00000000000000000000000011111110";
B14<= "00000000000000000000000011111110";
B15<= "00000000000000000000000000000111";
B16<= "00000000000000000000000000000000";
B17<= "00000000000000000000000000000000";
B18<= "00000000000000000000000000000000";
B19<= "00000000000000000000000000000000";
B20<= "00000000000000000000000000000000";
B21<= "00000000000000000000000000000000";
B22<= "00000000000000000000000000000000";
B23<= "00000000000000000000000000000000";
B24<= "00000000000000000000000000000000";
B25<= "00000000000000000000000000000000";
B26<= "00000000000000000000000000000000";

process (x, y, x_en, y_en, draw_count)
begin
	if (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 32) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R1(to_integer(unsigned(draw_count)));
			G <= G1(to_integer(unsigned(draw_count)));
			B <= B1(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 33) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R2(to_integer(unsigned(draw_count)));
			G <= G2(to_integer(unsigned(draw_count)));
			B <= B2(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 34) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R3(to_integer(unsigned(draw_count)));
			G <= G3(to_integer(unsigned(draw_count)));
			B <= B3(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 35) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R4(to_integer(unsigned(draw_count)));
			G <= G4(to_integer(unsigned(draw_count)));
			B <= B4(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 36) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R5(to_integer(unsigned(draw_count)));
			G <= G5(to_integer(unsigned(draw_count)));
			B <= B5(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 37) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R6(to_integer(unsigned(draw_count)));
			G <= G6(to_integer(unsigned(draw_count)));
			B <= B6(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 38) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R7(to_integer(unsigned(draw_count)));
			G <= G7(to_integer(unsigned(draw_count)));
			B <= B7(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 39) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R8(to_integer(unsigned(draw_count)));
			G <= G8(to_integer(unsigned(draw_count)));
			B <= B8(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 40) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R9(to_integer(unsigned(draw_count)));
			G <= G9(to_integer(unsigned(draw_count)));
			B <= B9(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 41) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R10(to_integer(unsigned(draw_count)));
			G <= G10(to_integer(unsigned(draw_count)));
			B <= B10(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 42) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R11(to_integer(unsigned(draw_count)));
			G <= G11(to_integer(unsigned(draw_count)));
			B <= B11(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 43) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R12(to_integer(unsigned(draw_count)));
			G <= G12(to_integer(unsigned(draw_count)));
			B <= B12(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 44) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R13(to_integer(unsigned(draw_count)));
			G <= G13(to_integer(unsigned(draw_count)));
			B <= B13(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 45) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R14(to_integer(unsigned(draw_count)));
			G <= G14(to_integer(unsigned(draw_count)));
			B <= B14(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 46) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R15(to_integer(unsigned(draw_count)));
			G <= G15(to_integer(unsigned(draw_count)));
			B <= B15(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 47) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R16(to_integer(unsigned(draw_count)));
			G <= G16(to_integer(unsigned(draw_count)));
			B <= B16(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 48) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R17(to_integer(unsigned(draw_count)));
			G <= G17(to_integer(unsigned(draw_count)));
			B <= B17(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 49) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R18(to_integer(unsigned(draw_count)));
			G <= G18(to_integer(unsigned(draw_count)));
			B <= B18(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 50) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R19(to_integer(unsigned(draw_count)));
			G <= G19(to_integer(unsigned(draw_count)));
			B <= B19(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 51) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R20(to_integer(unsigned(draw_count)));
			G <= G20(to_integer(unsigned(draw_count)));
			B <= B20(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 52) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R21(to_integer(unsigned(draw_count)));
			G <= G21(to_integer(unsigned(draw_count)));
			B <= B21(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 53) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R22(to_integer(unsigned(draw_count)));
			G <= G22(to_integer(unsigned(draw_count)));
			B <= B22(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 54) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R23(to_integer(unsigned(draw_count)));
			G <= G23(to_integer(unsigned(draw_count)));
			B <= B23(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 55) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R24(to_integer(unsigned(draw_count)));
			G <= G24(to_integer(unsigned(draw_count)));
			B <= B24(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 56) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R25(to_integer(unsigned(draw_count)));
			G <= G25(to_integer(unsigned(draw_count)));
			B <= B25(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	elsif (to_integer(unsigned(y)) = to_integer(unsigned(y_en)) + 57) then	
		if (to_integer(unsigned(x)) >= to_integer(unsigned(x_en)) + 69 and 
		to_integer(unsigned(x)) <= to_integer(unsigned(x_en)) + 100) then
			enable <= '1';
			R <= R26(to_integer(unsigned(draw_count)));
			G <= G26(to_integer(unsigned(draw_count)));
			B <= B26(to_integer(unsigned(draw_count)));
		else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
		end if;
	else
			enable <= '0';
			R <= '0';
			G <= '0';
			B <= '0';
	end if;
end process;	

end behaviour;

