library IEEE;
use IEEE.std_logic_1164.ALL;

architecture behaviour of draw_title is
begin

r <= gameover;
g <= '0';
b <= menu;

end behaviour;

