configuration draw_counter_behaviour_cfg of draw_counter is
   for behaviour
   end for;
end draw_counter_behaviour_cfg;
