
library ieee;
use ieee.std_logic_1164.all;
--library tcb018gbwp7t;
--use tcb018gbwp7t.all;

architecture synthesised of display is

  component INVD4BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component ND2D4BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INR3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component NR4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component OR4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component OR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component OAI211D1BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component AOI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component OAI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component AOI211XD0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component AN4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component IND4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component AOI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component IOA21D1BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component AO21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component OA31D1BWP7T
    port(A1, A2, A3, B : in std_logic; Z : out std_logic);
  end component;

  component OAI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OAI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component OAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component NR3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component CKAN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component NR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INVD0BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component MOAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component IAO21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component AOI32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component ND3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component AN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component CKND1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component IND3D1BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component ND4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component INVD1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component AOI211D1BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component OA22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component INR2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component AOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2XD0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component IND2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component OR3D1BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component INR4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component AN3D1BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component AN2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component INR2XD0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component OA21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component MAOI222D1BWP7T
    port(A, B, C : in std_logic; ZN : out std_logic);
  end component;

  component AN3D0BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component MAOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component CKND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component CKND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component XNR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component IIND4D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component CKXOR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component DFCNQD1BWP7T
    port(CDN, CP, D : in std_logic; Q : out std_logic);
  end component;

  component AO31D1BWP7T
    port(A1, A2, A3, B : in std_logic; Z : out std_logic);
  end component;

  component AO211D0BWP7T
    port(A1, A2, B, C : in std_logic; Z : out std_logic);
  end component;

  component INR2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component IND2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component AO221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component OAI32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component AOI211D0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component OA211D0BWP7T
    port(A1, A2, B, C : in std_logic; Z : out std_logic);
  end component;

  component DFQD1BWP7T
    port(CP, D : in std_logic; Q : out std_logic);
  end component;

  component OAI32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component DFD1BWP7T
    port(CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component AO22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component DFXQD1BWP7T
    port(CP, DA, DB, SA : in std_logic; Q : out std_logic);
  end component;

  signal x : std_logic_vector(8 downto 0);
  signal y : std_logic_vector(9 downto 0);
  signal draw_count4 : std_logic_vector(4 downto 0);
  signal draw_count2 : std_logic_vector(4 downto 0);
  signal draw_count3 : std_logic_vector(4 downto 0);
  signal draw_count5 : std_logic_vector(4 downto 0);
  signal draw_count6 : std_logic_vector(4 downto 0);
  signal draw_count7 : std_logic_vector(4 downto 0);
  signal draw_count8 : std_logic_vector(4 downto 0);
  signal draw_count10 : std_logic_vector(4 downto 0);
  signal draw_count9 : std_logic_vector(4 downto 0);
  signal draw_count1 : std_logic_vector(4 downto 0);
  signal UNCONNECTED, UNCONNECTED0, b1, b2, b3 : std_logic;
  signal b4, b5, b6, b7, b8 : std_logic;
  signal b9, b10, enable1, enable2, enable3 : std_logic;
  signal enable4, enable5, enable6, enable7, enable8 : std_logic;
  signal enable9, enable10, g1, g2, g3 : std_logic;
  signal g4, g5, g6, g7, g8 : std_logic;
  signal g9, g10, l01_n_0, l01_n_1, l01_n_2 : std_logic;
  signal l01_n_3, l01_n_4, l01_n_5, l01_n_6, l01_n_7 : std_logic;
  signal l01_n_8, l01_n_9, l01_n_10, l01_n_11, l01_n_12 : std_logic;
  signal l01_n_13, l01_n_14, l01_n_15, l01_n_16, l01_n_17 : std_logic;
  signal l01_n_18, l01_n_19, l01_n_20, l01_n_21, l01_n_22 : std_logic;
  signal l01_n_23, l01_n_24, l01_n_25, l01_n_26, l01_n_27 : std_logic;
  signal l01_n_28, l01_n_29, l01_n_30, l01_n_31, l02_n_0 : std_logic;
  signal l02_n_1, l02_n_3, l02_n_4, l02_n_5, l02_n_6 : std_logic;
  signal l02_n_7, l02_n_8, l02_n_9, l02_n_10, l02_n_11 : std_logic;
  signal l02_n_12, l02_n_13, l02_n_14, l02_n_15, l02_n_16 : std_logic;
  signal l02_n_17, l02_n_18, l02_n_19, l02_n_20, l02_n_21 : std_logic;
  signal l02_n_22, l02_n_23, l02_n_24, l02_n_25, l02_n_26 : std_logic;
  signal l02_n_27, l02_n_28, l02_n_29, l02_n_30, l02_n_31 : std_logic;
  signal l02_n_32, l02_n_33, l02_n_34, l02_n_35, l02_n_36 : std_logic;
  signal l02_n_37, l02_n_38, l02_n_39, l03_n_0, l03_n_1 : std_logic;
  signal l03_n_2, l03_n_3, l03_n_4, l03_n_5, l03_n_6 : std_logic;
  signal l03_n_7, l03_n_9, l03_n_11, l03_n_33, l03_vold : std_logic;
  signal l06_n_0, l06_n_1, l06_n_2, l06_n_3, l06_n_4 : std_logic;
  signal l06_n_5, l06_n_6, l06_n_7, l06_n_8, l06_n_9 : std_logic;
  signal l06_n_10, l06_n_11, l06_n_12, l06_n_13, l06_n_14 : std_logic;
  signal l06_n_15, l06_n_16, l06_n_17, l06_n_18, l06_n_19 : std_logic;
  signal l06_n_20, l06_n_21, l06_n_22, l06_n_23, l06_n_24 : std_logic;
  signal l06_n_25, l06_n_26, l06_n_27, l06_n_28, l06_n_29 : std_logic;
  signal l06_n_30, l06_n_31, l06_n_32, l06_n_33, l06_n_34 : std_logic;
  signal l06_n_35, l06_n_36, l06_n_37, l06_n_38, l06_n_39 : std_logic;
  signal l06_n_41, l06_n_42, l06_n_43, l06_n_44, l06_n_45 : std_logic;
  signal l06_n_46, l06_n_47, l06_n_48, l06_n_49, l06_n_50 : std_logic;
  signal l06_n_51, l06_n_52, l06_n_53, l06_n_54, l06_n_56 : std_logic;
  signal l06_n_57, l06_n_58, l06_n_59, l06_n_60, l06_n_61 : std_logic;
  signal l06_n_62, l06_n_63, l06_n_64, l06_n_65, l06_n_66 : std_logic;
  signal l06_n_67, l06_n_68, l06_n_69, l06_n_70, l06_n_71 : std_logic;
  signal l06_n_72, l06_n_73, l06_n_74, l06_n_75, l06_n_76 : std_logic;
  signal l06_n_77, l06_n_78, l06_n_79, l06_n_80, l06_n_81 : std_logic;
  signal l06_n_82, l06_n_83, l06_n_84, l06_n_85, l06_n_86 : std_logic;
  signal l06_n_87, l06_n_88, l06_n_89, l06_n_90, l06_n_91 : std_logic;
  signal l06_n_92, l06_n_93, l06_n_95, l06_n_96, l06_n_97 : std_logic;
  signal l06_n_98, l06_n_99, l06_n_100, l06_n_101, l06_n_104 : std_logic;
  signal l06_n_105, l06_n_106, l06_n_107, l06_n_108, l06_n_109 : std_logic;
  signal l06_n_110, l06_n_111, l06_n_112, l06_n_113, l06_n_114 : std_logic;
  signal l06_n_115, l06_n_116, l06_n_117, l06_n_118, l06_n_119 : std_logic;
  signal l06_n_120, l06_n_121, l06_n_122, l06_n_123, l06_n_124 : std_logic;
  signal l06_n_125, l06_n_126, l06_n_127, l06_n_128, l06_n_129 : std_logic;
  signal l06_n_130, l06_n_131, l06_n_132, l06_n_133, l06_n_134 : std_logic;
  signal l06_n_135, l06_n_136, l06_n_137, l06_n_138, l06_n_139 : std_logic;
  signal l06_n_140, l06_n_141, l06_n_142, l06_n_143, l06_n_144 : std_logic;
  signal l06_n_145, l06_n_146, l06_n_147, l06_n_148, l06_n_149 : std_logic;
  signal l06_n_150, l06_n_151, l06_n_152, l06_n_153, l06_n_154 : std_logic;
  signal l06_n_155, l06_n_156, l06_n_157, l06_n_158, l06_n_159 : std_logic;
  signal l06_n_160, l06_n_161, l06_n_162, l06_n_163, l06_n_164 : std_logic;
  signal l06_n_165, l06_n_166, l06_n_167, l06_n_168, l06_n_169 : std_logic;
  signal l06_n_170, l06_n_171, l06_n_172, l06_n_173, l06_n_174 : std_logic;
  signal l06_n_175, l06_n_176, l06_n_177, l06_n_178, l06_n_179 : std_logic;
  signal l06_n_180, l06_n_181, l06_n_182, l06_n_183, l06_n_184 : std_logic;
  signal l06_n_185, l06_n_186, l06_n_187, l06_n_188, l06_n_189 : std_logic;
  signal l06_n_190, l06_n_191, l06_n_192, l06_n_193, l06_n_194 : std_logic;
  signal l06_n_195, l06_n_196, l06_n_197, l06_n_198, l06_n_199 : std_logic;
  signal l06_n_200, l06_n_201, l06_n_202, l06_n_203, l06_n_204 : std_logic;
  signal l06_n_205, l06_n_206, l06_n_207, l06_n_208, l06_n_209 : std_logic;
  signal l06_n_210, l06_n_211, l06_n_212, l06_n_213, l06_n_214 : std_logic;
  signal l06_n_215, l06_n_216, l06_n_217, l06_n_218, l06_n_219 : std_logic;
  signal l06_n_220, l06_n_221, l06_n_222, l06_n_223, l06_n_224 : std_logic;
  signal l06_n_225, l06_n_226, l06_n_227, l06_n_228, l06_n_229 : std_logic;
  signal l06_n_230, l06_n_231, l06_n_232, l06_n_233, l06_n_234 : std_logic;
  signal l06_n_235, l06_n_236, l06_n_237, l06_n_238, l06_n_239 : std_logic;
  signal l06_n_240, l06_n_241, l06_n_242, l06_n_243, l06_n_244 : std_logic;
  signal l06_n_245, l06_n_246, l06_n_247, l06_n_248, l06_n_249 : std_logic;
  signal l06_n_250, l06_n_251, l06_n_252, l06_n_253, l06_n_254 : std_logic;
  signal l06_n_255, l06_n_256, l06_n_257, l06_n_258, l06_n_259 : std_logic;
  signal l06_n_260, l06_n_261, l06_n_262, l06_n_263, l06_n_264 : std_logic;
  signal l06_n_265, l06_n_266, l06_n_267, l06_n_268, l06_n_269 : std_logic;
  signal l06_n_270, l06_n_271, l06_n_272, l06_n_273, l06_n_274 : std_logic;
  signal l06_n_275, l06_n_276, l06_n_277, l06_n_278, l06_n_279 : std_logic;
  signal l06_n_280, l06_n_281, l06_n_282, l06_n_283, l06_n_284 : std_logic;
  signal l06_n_285, l06_n_286, l06_n_287, l06_n_288, l06_n_289 : std_logic;
  signal l06_n_290, l06_n_291, l06_n_292, l06_n_293, l06_n_294 : std_logic;
  signal l06_n_295, l06_n_296, l06_n_297, l06_n_298, l06_n_299 : std_logic;
  signal l06_n_300, l06_n_301, l06_n_302, l06_n_303, l06_n_304 : std_logic;
  signal l06_n_305, l06_n_306, l06_n_307, l06_n_308, l06_n_309 : std_logic;
  signal l06_n_311, l06_n_312, l06_n_313, l06_n_314, l06_n_315 : std_logic;
  signal l06_n_316, l06_n_317, l06_n_318, l06_n_319, l06_n_320 : std_logic;
  signal l06_n_321, l06_n_322, l06_n_323, l06_n_324, l06_n_325 : std_logic;
  signal l06_n_371, l06_n_372, l041_n_0, l041_n_1, l041_n_2 : std_logic;
  signal l041_n_3, l041_n_4, l041_n_5, l041_n_6, l042_n_0 : std_logic;
  signal l042_n_1, l042_n_2, l042_n_3, l042_n_4, l042_n_5 : std_logic;
  signal l042_n_6, l043_n_0, l043_n_1, l043_n_2, l043_n_3 : std_logic;
  signal l043_n_4, l043_n_5, l043_n_6, l044_n_0, l044_n_1 : std_logic;
  signal l044_n_2, l044_n_3, l044_n_4, l044_n_5, l044_n_6 : std_logic;
  signal l044_n_7, l044_n_8, l044_n_9, l044_n_10, l044_n_11 : std_logic;
  signal l044_n_12, l045_n_0, l045_n_1, l045_n_2, l045_n_3 : std_logic;
  signal l045_n_4, l045_n_5, l045_n_6, l045_n_7, l045_n_8 : std_logic;
  signal l045_n_9, l045_n_10, l045_n_11, l045_n_12, l046_n_0 : std_logic;
  signal l046_n_1, l046_n_2, l046_n_3, l046_n_4, l046_n_5 : std_logic;
  signal l046_n_6, l046_n_7, l046_n_8, l046_n_9, l046_n_10 : std_logic;
  signal l046_n_11, l046_n_12, l047_n_0, l047_n_1, l047_n_2 : std_logic;
  signal l047_n_3, l047_n_4, l047_n_5, l047_n_6, l047_n_7 : std_logic;
  signal l047_n_8, l047_n_9, l047_n_10, l047_n_11, l047_n_12 : std_logic;
  signal l048_n_0, l048_n_1, l048_n_2, l048_n_3, l048_n_4 : std_logic;
  signal l048_n_5, l048_n_6, l048_n_7, l048_n_8, l048_n_9 : std_logic;
  signal l048_n_10, l048_n_11, l048_n_12, l049_n_0, l049_n_1 : std_logic;
  signal l049_n_2, l049_n_3, l049_n_4, l049_n_5, l049_n_6 : std_logic;
  signal l049_n_7, l049_n_8, l049_n_9, l049_n_10, l049_n_11 : std_logic;
  signal l049_n_12, l051_n_0, l051_n_1, l051_n_2, l051_n_3 : std_logic;
  signal l051_n_4, l051_n_5, l051_n_6, l051_n_7, l051_n_8 : std_logic;
  signal l051_n_9, l051_n_10, l051_n_11, l051_n_12, l051_n_13 : std_logic;
  signal l051_n_14, l051_n_15, l051_n_16, l051_n_17, l051_n_18 : std_logic;
  signal l051_n_19, l051_n_20, l051_n_21, l051_n_22, l051_n_23 : std_logic;
  signal l051_n_24, l051_n_25, l051_n_26, l051_n_27, l051_n_28 : std_logic;
  signal l051_n_29, l051_n_30, l051_n_31, l051_n_32, l051_n_33 : std_logic;
  signal l051_n_34, l051_n_35, l051_n_36, l051_n_37, l051_n_38 : std_logic;
  signal l051_n_39, l051_n_40, l051_n_41, l051_n_42, l051_n_43 : std_logic;
  signal l051_n_44, l051_n_45, l051_n_46, l051_n_47, l051_n_48 : std_logic;
  signal l051_n_49, l051_n_50, l051_n_51, l051_n_52, l051_n_53 : std_logic;
  signal l051_n_54, l051_n_55, l051_n_56, l051_n_57, l051_n_58 : std_logic;
  signal l051_n_59, l051_n_60, l051_n_61, l051_n_62, l051_n_63 : std_logic;
  signal l051_n_64, l051_n_65, l051_n_66, l051_n_67, l051_n_68 : std_logic;
  signal l051_n_69, l051_n_70, l051_n_71, l051_n_72, l051_n_73 : std_logic;
  signal l051_n_74, l051_n_75, l051_n_76, l051_n_77, l051_n_78 : std_logic;
  signal l051_n_79, l051_n_80, l051_n_82, l051_n_83, l052_n_0 : std_logic;
  signal l052_n_1, l052_n_2, l052_n_3, l052_n_4, l052_n_5 : std_logic;
  signal l052_n_6, l052_n_7, l052_n_8, l052_n_9, l052_n_10 : std_logic;
  signal l052_n_11, l052_n_12, l052_n_13, l052_n_14, l052_n_15 : std_logic;
  signal l052_n_16, l052_n_17, l052_n_18, l052_n_19, l052_n_20 : std_logic;
  signal l052_n_21, l052_n_22, l052_n_23, l052_n_24, l052_n_25 : std_logic;
  signal l052_n_26, l052_n_27, l052_n_28, l052_n_29, l052_n_30 : std_logic;
  signal l052_n_31, l052_n_32, l052_n_33, l052_n_34, l052_n_35 : std_logic;
  signal l052_n_36, l052_n_37, l052_n_38, l052_n_39, l052_n_40 : std_logic;
  signal l052_n_41, l052_n_42, l052_n_43, l052_n_44, l052_n_45 : std_logic;
  signal l052_n_46, l052_n_47, l052_n_48, l052_n_49, l052_n_50 : std_logic;
  signal l052_n_51, l052_n_52, l052_n_53, l052_n_54, l052_n_55 : std_logic;
  signal l052_n_56, l052_n_57, l052_n_58, l052_n_59, l052_n_60 : std_logic;
  signal l052_n_61, l052_n_62, l052_n_63, l052_n_64, l052_n_65 : std_logic;
  signal l052_n_66, l052_n_67, l052_n_68, l052_n_69, l052_n_70 : std_logic;
  signal l052_n_71, l052_n_72, l052_n_73, l052_n_74, l052_n_75 : std_logic;
  signal l052_n_76, l052_n_77, l052_n_78, l052_n_79, l052_n_80 : std_logic;
  signal l052_n_82, l052_n_83, l053_n_0, l053_n_1, l053_n_2 : std_logic;
  signal l053_n_3, l053_n_4, l053_n_5, l053_n_6, l053_n_7 : std_logic;
  signal l053_n_8, l053_n_9, l053_n_10, l053_n_11, l053_n_12 : std_logic;
  signal l053_n_13, l053_n_14, l053_n_15, l053_n_16, l053_n_17 : std_logic;
  signal l053_n_18, l053_n_19, l053_n_20, l053_n_21, l053_n_22 : std_logic;
  signal l053_n_23, l053_n_24, l053_n_25, l053_n_26, l053_n_27 : std_logic;
  signal l053_n_28, l053_n_29, l053_n_30, l053_n_31, l053_n_32 : std_logic;
  signal l053_n_33, l053_n_34, l053_n_35, l053_n_36, l053_n_37 : std_logic;
  signal l053_n_38, l053_n_39, l053_n_40, l053_n_41, l053_n_42 : std_logic;
  signal l053_n_43, l053_n_44, l053_n_45, l053_n_46, l053_n_47 : std_logic;
  signal l053_n_48, l053_n_49, l053_n_50, l053_n_51, l053_n_52 : std_logic;
  signal l053_n_53, l053_n_54, l053_n_55, l053_n_56, l053_n_57 : std_logic;
  signal l053_n_58, l053_n_59, l053_n_60, l053_n_61, l053_n_62 : std_logic;
  signal l053_n_63, l053_n_64, l053_n_65, l053_n_66, l053_n_67 : std_logic;
  signal l053_n_68, l053_n_69, l053_n_70, l053_n_71, l053_n_72 : std_logic;
  signal l053_n_73, l053_n_74, l053_n_75, l053_n_76, l053_n_77 : std_logic;
  signal l053_n_78, l053_n_79, l053_n_80, l053_n_82, l053_n_83 : std_logic;
  signal l071_n_0, l071_n_1, l071_n_2, l071_n_3, l071_n_4 : std_logic;
  signal l071_n_5, l071_n_6, l071_n_7, l071_n_8, l071_n_9 : std_logic;
  signal l071_n_10, l071_n_11, l071_n_12, l071_n_13, l071_n_14 : std_logic;
  signal l071_n_15, l071_n_16, l071_n_17, l071_n_18, l071_n_19 : std_logic;
  signal l071_n_20, l071_n_21, l071_n_22, l071_n_23, l071_n_24 : std_logic;
  signal l071_n_25, l071_n_26, l071_n_27, l071_n_28, l071_n_29 : std_logic;
  signal l071_n_30, l071_n_31, l071_n_32, l071_n_33, l071_n_34 : std_logic;
  signal l071_n_35, l071_n_36, l071_n_37, l071_n_38, l071_n_39 : std_logic;
  signal l071_n_40, l071_n_41, l071_n_42, l071_n_43, l071_n_44 : std_logic;
  signal l071_n_45, l071_n_46, l071_n_47, l071_n_48, l071_n_49 : std_logic;
  signal l071_n_50, l071_n_51, l071_n_52, l071_n_53, l071_n_54 : std_logic;
  signal l071_n_55, l071_n_56, l071_n_57, l071_n_58, l071_n_59 : std_logic;
  signal l071_n_60, l071_n_61, l071_n_62, l071_n_63, l071_n_64 : std_logic;
  signal l071_n_65, l071_n_66, l071_n_67, l071_n_68, l071_n_69 : std_logic;
  signal l071_n_70, l071_n_71, l071_n_72, l071_n_73, l071_n_74 : std_logic;
  signal l071_n_75, l071_n_76, l071_n_77, l071_n_78, l071_n_79 : std_logic;
  signal l071_n_80, l071_n_81, l071_n_82, l071_n_83, l071_n_84 : std_logic;
  signal l071_n_85, l071_n_86, l071_n_87, l071_n_88, l071_n_89 : std_logic;
  signal l071_n_90, l071_n_91, l071_n_92, l071_n_93, l071_n_94 : std_logic;
  signal l071_n_95, l071_n_96, l071_n_97, l071_n_98, l071_n_99 : std_logic;
  signal l071_n_100, l071_n_101, l071_n_102, l071_n_103, l071_n_104 : std_logic;
  signal l071_n_105, l071_n_106, l071_n_107, l071_n_108, l071_n_109 : std_logic;
  signal l071_n_110, l071_n_111, l071_n_112, l071_n_113, l071_n_114 : std_logic;
  signal l071_n_115, l071_n_116, l071_n_117, l071_n_118, l071_n_119 : std_logic;
  signal l071_n_120, l071_n_121, l071_n_122, l071_n_123, l071_n_124 : std_logic;
  signal l071_n_125, l071_n_126, l071_n_127, l071_n_128, l071_n_129 : std_logic;
  signal l071_n_130, l071_n_131, l071_n_132, l071_n_133, l071_n_134 : std_logic;
  signal l071_n_135, l071_n_136, l071_n_137, l071_n_138, l071_n_139 : std_logic;
  signal l071_n_140, l071_n_141, l071_n_142, l071_n_143, l071_n_144 : std_logic;
  signal l071_n_145, l071_n_146, l071_n_147, l071_n_148, l071_n_149 : std_logic;
  signal l071_n_150, l071_n_151, l071_n_152, l071_n_153, l071_n_154 : std_logic;
  signal l071_n_155, l071_n_156, l071_n_157, l071_n_158, l071_n_159 : std_logic;
  signal l071_n_160, l071_n_161, l071_n_162, l071_n_163, l071_n_164 : std_logic;
  signal l071_n_165, l071_n_166, l071_n_167, l071_n_168, l071_n_169 : std_logic;
  signal l071_n_170, l071_n_171, l071_n_172, l071_n_173, l071_n_174 : std_logic;
  signal l071_n_175, l071_n_176, l071_n_177, l071_n_178, l071_n_179 : std_logic;
  signal l071_n_180, l071_n_181, l071_n_182, l071_n_183, l071_n_184 : std_logic;
  signal l071_n_185, l071_n_186, l071_n_187, l071_n_188, l071_n_189 : std_logic;
  signal l071_n_190, l071_n_191, l071_n_192, l071_n_193, l071_n_194 : std_logic;
  signal l071_n_195, l071_n_196, l071_n_197, l071_n_198, l071_n_199 : std_logic;
  signal l071_n_200, l071_n_201, l071_n_202, l071_n_203, l071_n_204 : std_logic;
  signal l071_n_205, l071_n_206, l071_n_207, l071_n_208, l071_n_209 : std_logic;
  signal l071_n_210, l071_n_211, l071_n_212, l071_n_213, l071_n_214 : std_logic;
  signal l071_n_215, l071_n_216, l071_n_217, l071_n_218, l071_n_219 : std_logic;
  signal l071_n_220, l071_n_221, l071_n_222, l071_n_223, l071_n_224 : std_logic;
  signal l071_n_225, l071_n_226, l071_n_227, l071_n_228, l071_n_229 : std_logic;
  signal l071_n_230, l071_n_231, l071_n_232, l071_n_233, l071_n_234 : std_logic;
  signal l071_n_235, l071_n_236, l071_n_237, l071_n_239, l071_n_241 : std_logic;
  signal l071_n_242, l071_n_243, l071_n_245, l071_n_246, l072_n_0 : std_logic;
  signal l072_n_1, l072_n_2, l072_n_3, l072_n_4, l072_n_5 : std_logic;
  signal l072_n_6, l072_n_7, l072_n_8, l072_n_9, l072_n_10 : std_logic;
  signal l072_n_11, l072_n_12, l072_n_13, l072_n_14, l072_n_15 : std_logic;
  signal l072_n_16, l072_n_17, l072_n_18, l072_n_19, l072_n_20 : std_logic;
  signal l072_n_21, l072_n_22, l072_n_23, l072_n_24, l072_n_25 : std_logic;
  signal l072_n_26, l072_n_27, l072_n_28, l072_n_29, l072_n_30 : std_logic;
  signal l072_n_31, l072_n_32, l072_n_33, l072_n_34, l072_n_35 : std_logic;
  signal l072_n_36, l072_n_37, l072_n_38, l072_n_39, l072_n_40 : std_logic;
  signal l072_n_41, l072_n_42, l072_n_43, l072_n_44, l072_n_45 : std_logic;
  signal l072_n_46, l072_n_47, l072_n_48, l072_n_49, l072_n_50 : std_logic;
  signal l072_n_51, l072_n_52, l072_n_53, l072_n_54, l072_n_55 : std_logic;
  signal l072_n_56, l072_n_57, l072_n_58, l072_n_59, l072_n_60 : std_logic;
  signal l072_n_61, l072_n_62, l072_n_63, l072_n_64, l072_n_65 : std_logic;
  signal l072_n_66, l072_n_67, l072_n_68, l072_n_69, l072_n_70 : std_logic;
  signal l072_n_71, l072_n_72, l072_n_73, l072_n_74, l072_n_75 : std_logic;
  signal l072_n_76, l072_n_77, l072_n_78, l072_n_79, l072_n_80 : std_logic;
  signal l072_n_81, l072_n_82, l072_n_83, l072_n_84, l072_n_85 : std_logic;
  signal l072_n_86, l072_n_87, l072_n_88, l072_n_89, l072_n_90 : std_logic;
  signal l072_n_91, l072_n_92, l072_n_93, l072_n_94, l072_n_95 : std_logic;
  signal l072_n_96, l072_n_97, l072_n_98, l072_n_99, l072_n_100 : std_logic;
  signal l072_n_101, l072_n_102, l072_n_103, l072_n_104, l072_n_105 : std_logic;
  signal l072_n_106, l072_n_107, l072_n_108, l072_n_109, l072_n_110 : std_logic;
  signal l072_n_111, l072_n_112, l072_n_113, l072_n_114, l072_n_115 : std_logic;
  signal l072_n_116, l072_n_117, l072_n_118, l072_n_119, l072_n_120 : std_logic;
  signal l072_n_121, l072_n_122, l072_n_123, l072_n_124, l072_n_125 : std_logic;
  signal l072_n_126, l072_n_127, l072_n_128, l072_n_129, l072_n_130 : std_logic;
  signal l072_n_131, l072_n_132, l072_n_133, l072_n_134, l072_n_135 : std_logic;
  signal l072_n_136, l072_n_137, l072_n_138, l072_n_139, l072_n_140 : std_logic;
  signal l072_n_141, l072_n_142, l072_n_143, l072_n_144, l072_n_145 : std_logic;
  signal l072_n_146, l072_n_147, l072_n_148, l072_n_149, l072_n_150 : std_logic;
  signal l072_n_151, l072_n_152, l072_n_153, l072_n_154, l072_n_155 : std_logic;
  signal l072_n_156, l072_n_157, l072_n_158, l072_n_159, l072_n_160 : std_logic;
  signal l072_n_161, l072_n_162, l072_n_163, l072_n_164, l072_n_165 : std_logic;
  signal l072_n_166, l072_n_167, l072_n_168, l072_n_169, l072_n_170 : std_logic;
  signal l072_n_171, l072_n_172, l072_n_173, l072_n_174, l072_n_175 : std_logic;
  signal l072_n_176, l072_n_177, l072_n_178, l072_n_179, l072_n_180 : std_logic;
  signal l072_n_181, l072_n_182, l072_n_183, l072_n_184, l072_n_185 : std_logic;
  signal l072_n_186, l072_n_187, l072_n_188, l072_n_189, l072_n_190 : std_logic;
  signal l072_n_191, l072_n_192, l072_n_193, l072_n_194, l072_n_195 : std_logic;
  signal l072_n_196, l072_n_197, l072_n_198, l072_n_199, l072_n_200 : std_logic;
  signal l072_n_201, l072_n_202, l072_n_203, l072_n_204, l072_n_205 : std_logic;
  signal l072_n_206, l072_n_207, l072_n_208, l072_n_209, l072_n_210 : std_logic;
  signal l072_n_211, l072_n_212, l072_n_213, l072_n_214, l072_n_215 : std_logic;
  signal l072_n_216, l072_n_217, l072_n_218, l072_n_219, l072_n_220 : std_logic;
  signal l072_n_221, l072_n_222, l072_n_223, l072_n_224, l072_n_225 : std_logic;
  signal l072_n_226, l072_n_227, l072_n_228, l072_n_229, l072_n_230 : std_logic;
  signal l072_n_231, l072_n_232, l072_n_233, l072_n_234, l072_n_235 : std_logic;
  signal l072_n_236, l072_n_237, l072_n_239, l072_n_241, l072_n_242 : std_logic;
  signal l072_n_243, l072_n_245, l072_n_246, l073_n_0, l073_n_1 : std_logic;
  signal l073_n_2, l073_n_3, l073_n_4, l073_n_5, l073_n_6 : std_logic;
  signal l073_n_7, l073_n_8, l073_n_9, l073_n_10, l073_n_11 : std_logic;
  signal l073_n_12, l073_n_13, l073_n_14, l073_n_15, l073_n_16 : std_logic;
  signal l073_n_17, l073_n_18, l073_n_19, l073_n_20, l073_n_21 : std_logic;
  signal l073_n_22, l073_n_23, l073_n_24, l073_n_25, l073_n_26 : std_logic;
  signal l073_n_27, l073_n_28, l073_n_29, l073_n_30, l073_n_31 : std_logic;
  signal l073_n_32, l073_n_33, l073_n_34, l073_n_35, l073_n_36 : std_logic;
  signal l073_n_37, l073_n_38, l073_n_39, l073_n_40, l073_n_41 : std_logic;
  signal l073_n_42, l073_n_43, l073_n_44, l073_n_45, l073_n_46 : std_logic;
  signal l073_n_47, l073_n_48, l073_n_49, l073_n_50, l073_n_51 : std_logic;
  signal l073_n_52, l073_n_53, l073_n_54, l073_n_55, l073_n_56 : std_logic;
  signal l073_n_57, l073_n_58, l073_n_59, l073_n_60, l073_n_61 : std_logic;
  signal l073_n_62, l073_n_63, l073_n_64, l073_n_65, l073_n_66 : std_logic;
  signal l073_n_67, l073_n_68, l073_n_69, l073_n_70, l073_n_71 : std_logic;
  signal l073_n_72, l073_n_73, l073_n_74, l073_n_75, l073_n_76 : std_logic;
  signal l073_n_77, l073_n_78, l073_n_79, l073_n_80, l073_n_81 : std_logic;
  signal l073_n_82, l073_n_83, l073_n_84, l073_n_85, l073_n_86 : std_logic;
  signal l073_n_87, l073_n_88, l073_n_89, l073_n_90, l073_n_91 : std_logic;
  signal l073_n_92, l073_n_93, l073_n_94, l073_n_95, l073_n_96 : std_logic;
  signal l073_n_97, l073_n_98, l073_n_99, l073_n_100, l073_n_101 : std_logic;
  signal l073_n_102, l073_n_103, l073_n_104, l073_n_105, l073_n_106 : std_logic;
  signal l073_n_107, l073_n_108, l073_n_109, l073_n_110, l073_n_111 : std_logic;
  signal l073_n_112, l073_n_113, l073_n_114, l073_n_115, l073_n_116 : std_logic;
  signal l073_n_117, l073_n_118, l073_n_119, l073_n_120, l073_n_121 : std_logic;
  signal l073_n_122, l073_n_123, l073_n_124, l073_n_125, l073_n_126 : std_logic;
  signal l073_n_127, l073_n_128, l073_n_129, l073_n_130, l073_n_131 : std_logic;
  signal l073_n_132, l073_n_133, l073_n_134, l073_n_135, l073_n_136 : std_logic;
  signal l073_n_137, l073_n_138, l073_n_139, l073_n_140, l073_n_141 : std_logic;
  signal l073_n_142, l073_n_143, l073_n_144, l073_n_145, l073_n_146 : std_logic;
  signal l073_n_147, l073_n_148, l073_n_149, l073_n_150, l073_n_151 : std_logic;
  signal l073_n_152, l073_n_153, l073_n_154, l073_n_155, l073_n_156 : std_logic;
  signal l073_n_157, l073_n_158, l073_n_159, l073_n_160, l073_n_161 : std_logic;
  signal l073_n_162, l073_n_163, l073_n_164, l073_n_165, l073_n_166 : std_logic;
  signal l073_n_167, l073_n_168, l073_n_169, l073_n_170, l073_n_171 : std_logic;
  signal l073_n_172, l073_n_173, l073_n_174, l073_n_175, l073_n_176 : std_logic;
  signal l073_n_177, l073_n_178, l073_n_179, l073_n_180, l073_n_181 : std_logic;
  signal l073_n_182, l073_n_183, l073_n_184, l073_n_185, l073_n_186 : std_logic;
  signal l073_n_187, l073_n_188, l073_n_189, l073_n_190, l073_n_191 : std_logic;
  signal l073_n_192, l073_n_193, l073_n_194, l073_n_195, l073_n_196 : std_logic;
  signal l073_n_197, l073_n_198, l073_n_199, l073_n_200, l073_n_201 : std_logic;
  signal l073_n_202, l073_n_203, l073_n_204, l073_n_205, l073_n_206 : std_logic;
  signal l073_n_207, l073_n_208, l073_n_209, l073_n_210, l073_n_211 : std_logic;
  signal l073_n_212, l073_n_213, l073_n_214, l073_n_215, l073_n_216 : std_logic;
  signal l073_n_217, l073_n_218, l073_n_219, l073_n_220, l073_n_221 : std_logic;
  signal l073_n_222, l073_n_223, l073_n_224, l073_n_225, l073_n_226 : std_logic;
  signal l073_n_227, l073_n_228, l073_n_229, l073_n_230, l073_n_231 : std_logic;
  signal l073_n_232, l073_n_233, l073_n_234, l073_n_235, l073_n_236 : std_logic;
  signal l073_n_237, l073_n_239, l073_n_241, l073_n_242, l073_n_243 : std_logic;
  signal l073_n_245, l073_n_246, l074_n_0, l074_n_1, l074_n_2 : std_logic;
  signal l074_n_3, l074_n_4, l074_n_5, l074_n_6, l074_n_7 : std_logic;
  signal l074_n_8, l074_n_9, l074_n_10, l074_n_11, l074_n_12 : std_logic;
  signal l074_n_13, l074_n_14, l074_n_15, l074_n_16, l074_n_17 : std_logic;
  signal l074_n_18, l074_n_19, l074_n_20, l074_n_21, l074_n_22 : std_logic;
  signal l074_n_23, l074_n_24, l074_n_25, l074_n_26, l074_n_27 : std_logic;
  signal l074_n_28, l074_n_29, l074_n_30, l074_n_31, l074_n_32 : std_logic;
  signal l074_n_33, l074_n_34, l074_n_35, l074_n_36, l074_n_37 : std_logic;
  signal l074_n_38, l074_n_39, l074_n_40, l074_n_41, l074_n_42 : std_logic;
  signal l074_n_43, l074_n_44, l074_n_45, l074_n_46, l074_n_47 : std_logic;
  signal l074_n_48, l074_n_49, l074_n_50, l074_n_51, l074_n_52 : std_logic;
  signal l074_n_53, l074_n_54, l074_n_55, l074_n_56, l074_n_57 : std_logic;
  signal l074_n_58, l074_n_59, l074_n_60, l074_n_61, l074_n_62 : std_logic;
  signal l074_n_63, l074_n_64, l074_n_65, l074_n_66, l074_n_67 : std_logic;
  signal l074_n_68, l074_n_69, l074_n_70, l074_n_71, l074_n_72 : std_logic;
  signal l074_n_73, l074_n_74, l074_n_75, l074_n_76, l074_n_77 : std_logic;
  signal l074_n_78, l074_n_79, l074_n_80, l074_n_81, l074_n_82 : std_logic;
  signal l074_n_83, l074_n_84, l074_n_85, l074_n_86, l074_n_87 : std_logic;
  signal l074_n_88, l074_n_89, l074_n_90, l074_n_91, l074_n_92 : std_logic;
  signal l074_n_93, l074_n_94, l074_n_95, l074_n_96, l074_n_97 : std_logic;
  signal l074_n_98, l074_n_99, l074_n_100, l074_n_101, l074_n_102 : std_logic;
  signal l074_n_103, l074_n_104, l074_n_105, l074_n_106, l074_n_107 : std_logic;
  signal l074_n_108, l074_n_109, l074_n_110, l074_n_111, l074_n_112 : std_logic;
  signal l074_n_113, l074_n_114, l074_n_115, l074_n_116, l074_n_117 : std_logic;
  signal l074_n_118, l074_n_119, l074_n_120, l074_n_121, l074_n_122 : std_logic;
  signal l074_n_123, l074_n_124, l074_n_125, l074_n_126, l074_n_127 : std_logic;
  signal l074_n_128, l074_n_129, l074_n_130, l074_n_131, l074_n_132 : std_logic;
  signal l074_n_133, l074_n_134, l074_n_135, l074_n_136, l074_n_137 : std_logic;
  signal l074_n_138, l074_n_139, l074_n_140, l074_n_141, l074_n_142 : std_logic;
  signal l074_n_143, l074_n_144, l074_n_145, l074_n_146, l074_n_147 : std_logic;
  signal l074_n_148, l074_n_149, l074_n_150, l074_n_151, l074_n_152 : std_logic;
  signal l074_n_153, l074_n_154, l074_n_155, l074_n_156, l074_n_157 : std_logic;
  signal l074_n_158, l074_n_159, l074_n_160, l074_n_161, l074_n_162 : std_logic;
  signal l074_n_163, l074_n_164, l074_n_165, l074_n_166, l074_n_167 : std_logic;
  signal l074_n_168, l074_n_169, l074_n_170, l074_n_171, l074_n_172 : std_logic;
  signal l074_n_173, l074_n_174, l074_n_175, l074_n_176, l074_n_177 : std_logic;
  signal l074_n_178, l074_n_179, l074_n_180, l074_n_181, l074_n_182 : std_logic;
  signal l074_n_183, l074_n_184, l074_n_185, l074_n_186, l074_n_187 : std_logic;
  signal l074_n_188, l074_n_189, l074_n_190, l074_n_191, l074_n_192 : std_logic;
  signal l074_n_193, l074_n_194, l074_n_195, l074_n_196, l074_n_197 : std_logic;
  signal l074_n_198, l074_n_199, l074_n_200, l074_n_201, l074_n_202 : std_logic;
  signal l074_n_203, l074_n_204, l074_n_205, l074_n_206, l074_n_207 : std_logic;
  signal l074_n_208, l074_n_209, l074_n_210, l074_n_211, l074_n_212 : std_logic;
  signal l074_n_213, l074_n_214, l074_n_215, l074_n_216, l074_n_217 : std_logic;
  signal l074_n_218, l074_n_219, l074_n_220, l074_n_221, l074_n_222 : std_logic;
  signal l074_n_223, l074_n_224, l074_n_225, l074_n_226, l074_n_227 : std_logic;
  signal l074_n_228, l074_n_229, l074_n_230, l074_n_231, l074_n_232 : std_logic;
  signal l074_n_233, l074_n_234, l074_n_235, l074_n_236, l074_n_238 : std_logic;
  signal l074_n_240, l074_n_241, l074_n_242, l074_n_244, l074_n_245 : std_logic;
  signal l075_n_0, l075_n_1, l075_n_2, l075_n_3, l075_n_4 : std_logic;
  signal l075_n_5, l075_n_6, l075_n_7, l075_n_8, l075_n_9 : std_logic;
  signal l075_n_10, l075_n_11, l075_n_12, l075_n_13, l075_n_14 : std_logic;
  signal l075_n_15, l075_n_16, l075_n_17, l075_n_18, l075_n_19 : std_logic;
  signal l075_n_20, l075_n_21, l075_n_22, l075_n_23, l075_n_24 : std_logic;
  signal l075_n_25, l075_n_26, l075_n_27, l075_n_28, l075_n_29 : std_logic;
  signal l075_n_30, l075_n_31, l075_n_32, l075_n_33, l075_n_34 : std_logic;
  signal l075_n_35, l075_n_36, l075_n_37, l075_n_38, l075_n_39 : std_logic;
  signal l075_n_40, l075_n_41, l075_n_42, l075_n_43, l075_n_44 : std_logic;
  signal l075_n_45, l075_n_46, l075_n_47, l075_n_48, l075_n_49 : std_logic;
  signal l075_n_50, l075_n_51, l075_n_52, l075_n_53, l075_n_54 : std_logic;
  signal l075_n_55, l075_n_56, l075_n_57, l075_n_58, l075_n_59 : std_logic;
  signal l075_n_60, l075_n_61, l075_n_62, l075_n_63, l075_n_64 : std_logic;
  signal l075_n_65, l075_n_66, l075_n_67, l075_n_68, l075_n_69 : std_logic;
  signal l075_n_70, l075_n_71, l075_n_72, l075_n_73, l075_n_74 : std_logic;
  signal l075_n_75, l075_n_76, l075_n_77, l075_n_78, l075_n_79 : std_logic;
  signal l075_n_80, l075_n_81, l075_n_82, l075_n_83, l075_n_84 : std_logic;
  signal l075_n_85, l075_n_86, l075_n_87, l075_n_88, l075_n_89 : std_logic;
  signal l075_n_90, l075_n_91, l075_n_92, l075_n_93, l075_n_94 : std_logic;
  signal l075_n_95, l075_n_96, l075_n_97, l075_n_98, l075_n_99 : std_logic;
  signal l075_n_100, l075_n_101, l075_n_102, l075_n_103, l075_n_104 : std_logic;
  signal l075_n_105, l075_n_106, l075_n_107, l075_n_108, l075_n_109 : std_logic;
  signal l075_n_110, l075_n_111, l075_n_112, l075_n_113, l075_n_114 : std_logic;
  signal l075_n_115, l075_n_116, l075_n_117, l075_n_118, l075_n_119 : std_logic;
  signal l075_n_120, l075_n_121, l075_n_122, l075_n_123, l075_n_124 : std_logic;
  signal l075_n_125, l075_n_126, l075_n_127, l075_n_128, l075_n_129 : std_logic;
  signal l075_n_130, l075_n_131, l075_n_132, l075_n_133, l075_n_134 : std_logic;
  signal l075_n_135, l075_n_136, l075_n_137, l075_n_138, l075_n_139 : std_logic;
  signal l075_n_140, l075_n_141, l075_n_142, l075_n_143, l075_n_144 : std_logic;
  signal l075_n_145, l075_n_146, l075_n_147, l075_n_148, l075_n_149 : std_logic;
  signal l075_n_150, l075_n_151, l075_n_152, l075_n_153, l075_n_154 : std_logic;
  signal l075_n_155, l075_n_156, l075_n_157, l075_n_158, l075_n_159 : std_logic;
  signal l075_n_160, l075_n_161, l075_n_162, l075_n_163, l075_n_164 : std_logic;
  signal l075_n_165, l075_n_166, l075_n_167, l075_n_168, l075_n_169 : std_logic;
  signal l075_n_170, l075_n_171, l075_n_172, l075_n_173, l075_n_174 : std_logic;
  signal l075_n_175, l075_n_176, l075_n_177, l075_n_178, l075_n_179 : std_logic;
  signal l075_n_180, l075_n_181, l075_n_182, l075_n_183, l075_n_184 : std_logic;
  signal l075_n_185, l075_n_186, l075_n_187, l075_n_188, l075_n_189 : std_logic;
  signal l075_n_190, l075_n_191, l075_n_192, l075_n_193, l075_n_194 : std_logic;
  signal l075_n_195, l075_n_196, l075_n_197, l075_n_198, l075_n_199 : std_logic;
  signal l075_n_200, l075_n_201, l075_n_202, l075_n_203, l075_n_204 : std_logic;
  signal l075_n_205, l075_n_206, l075_n_207, l075_n_208, l075_n_209 : std_logic;
  signal l075_n_210, l075_n_211, l075_n_212, l075_n_213, l075_n_214 : std_logic;
  signal l075_n_215, l075_n_216, l075_n_217, l075_n_218, l075_n_219 : std_logic;
  signal l075_n_220, l075_n_221, l075_n_222, l075_n_223, l075_n_224 : std_logic;
  signal l075_n_225, l075_n_226, l075_n_227, l075_n_228, l075_n_229 : std_logic;
  signal l075_n_230, l075_n_231, l075_n_232, l075_n_233, l075_n_234 : std_logic;
  signal l075_n_235, l075_n_236, l075_n_238, l075_n_240, l075_n_241 : std_logic;
  signal l075_n_242, l075_n_244, l075_n_245, l076_n_0, l076_n_1 : std_logic;
  signal l076_n_2, l076_n_3, l076_n_4, l076_n_5, l076_n_6 : std_logic;
  signal l076_n_7, l076_n_8, l076_n_9, l076_n_10, l076_n_11 : std_logic;
  signal l076_n_12, l076_n_13, l076_n_14, l076_n_15, l076_n_16 : std_logic;
  signal l076_n_17, l076_n_18, l076_n_19, l076_n_20, l076_n_21 : std_logic;
  signal l076_n_22, l076_n_23, l076_n_24, l076_n_25, l076_n_26 : std_logic;
  signal l076_n_27, l076_n_28, l076_n_29, l076_n_30, l076_n_31 : std_logic;
  signal l076_n_32, l076_n_33, l076_n_34, l076_n_35, l076_n_36 : std_logic;
  signal l076_n_37, l076_n_38, l076_n_39, l076_n_40, l076_n_41 : std_logic;
  signal l076_n_42, l076_n_43, l076_n_44, l076_n_45, l076_n_46 : std_logic;
  signal l076_n_47, l076_n_48, l076_n_49, l076_n_50, l076_n_51 : std_logic;
  signal l076_n_52, l076_n_53, l076_n_54, l076_n_55, l076_n_56 : std_logic;
  signal l076_n_57, l076_n_58, l076_n_59, l076_n_60, l076_n_61 : std_logic;
  signal l076_n_62, l076_n_63, l076_n_64, l076_n_65, l076_n_66 : std_logic;
  signal l076_n_67, l076_n_68, l076_n_69, l076_n_70, l076_n_71 : std_logic;
  signal l076_n_72, l076_n_73, l076_n_74, l076_n_75, l076_n_76 : std_logic;
  signal l076_n_77, l076_n_78, l076_n_79, l076_n_80, l076_n_81 : std_logic;
  signal l076_n_82, l076_n_83, l076_n_84, l076_n_85, l076_n_86 : std_logic;
  signal l076_n_87, l076_n_88, l076_n_89, l076_n_90, l076_n_91 : std_logic;
  signal l076_n_92, l076_n_93, l076_n_94, l076_n_95, l076_n_96 : std_logic;
  signal l076_n_97, l076_n_98, l076_n_99, l076_n_100, l076_n_101 : std_logic;
  signal l076_n_102, l076_n_103, l076_n_104, l076_n_105, l076_n_106 : std_logic;
  signal l076_n_107, l076_n_108, l076_n_109, l076_n_110, l076_n_111 : std_logic;
  signal l076_n_112, l076_n_113, l076_n_114, l076_n_115, l076_n_116 : std_logic;
  signal l076_n_117, l076_n_118, l076_n_119, l076_n_120, l076_n_121 : std_logic;
  signal l076_n_122, l076_n_123, l076_n_124, l076_n_125, l076_n_126 : std_logic;
  signal l076_n_127, l076_n_128, l076_n_129, l076_n_130, l076_n_131 : std_logic;
  signal l076_n_132, l076_n_133, l076_n_134, l076_n_135, l076_n_136 : std_logic;
  signal l076_n_137, l076_n_138, l076_n_139, l076_n_140, l076_n_141 : std_logic;
  signal l076_n_142, l076_n_143, l076_n_144, l076_n_145, l076_n_146 : std_logic;
  signal l076_n_147, l076_n_148, l076_n_149, l076_n_150, l076_n_151 : std_logic;
  signal l076_n_152, l076_n_153, l076_n_154, l076_n_155, l076_n_156 : std_logic;
  signal l076_n_157, l076_n_158, l076_n_159, l076_n_160, l076_n_161 : std_logic;
  signal l076_n_162, l076_n_163, l076_n_164, l076_n_165, l076_n_166 : std_logic;
  signal l076_n_167, l076_n_168, l076_n_169, l076_n_170, l076_n_171 : std_logic;
  signal l076_n_172, l076_n_173, l076_n_174, l076_n_175, l076_n_176 : std_logic;
  signal l076_n_177, l076_n_178, l076_n_179, l076_n_180, l076_n_181 : std_logic;
  signal l076_n_182, l076_n_183, l076_n_184, l076_n_185, l076_n_186 : std_logic;
  signal l076_n_187, l076_n_188, l076_n_189, l076_n_190, l076_n_191 : std_logic;
  signal l076_n_192, l076_n_193, l076_n_194, l076_n_195, l076_n_196 : std_logic;
  signal l076_n_197, l076_n_198, l076_n_199, l076_n_200, l076_n_201 : std_logic;
  signal l076_n_202, l076_n_203, l076_n_204, l076_n_205, l076_n_206 : std_logic;
  signal l076_n_207, l076_n_208, l076_n_209, l076_n_210, l076_n_211 : std_logic;
  signal l076_n_212, l076_n_213, l076_n_214, l076_n_215, l076_n_216 : std_logic;
  signal l076_n_217, l076_n_218, l076_n_219, l076_n_220, l076_n_221 : std_logic;
  signal l076_n_222, l076_n_223, l076_n_224, l076_n_225, l076_n_226 : std_logic;
  signal l076_n_227, l076_n_228, l076_n_229, l076_n_230, l076_n_231 : std_logic;
  signal l076_n_232, l076_n_233, l076_n_234, l076_n_235, l076_n_236 : std_logic;
  signal l076_n_238, l076_n_240, l076_n_241, l076_n_242, l076_n_244 : std_logic;
  signal l076_n_245, l0410_n_0, l0410_n_1, l0410_n_2, l0410_n_3 : std_logic;
  signal l0410_n_4, l0410_n_5, l0410_n_6, l0410_n_7, l0410_n_8 : std_logic;
  signal l0410_n_9, l0410_n_10, l0410_n_11, l0410_n_12, n_0 : std_logic;
  signal n_1, n_2, n_3, n_4, n_5 : std_logic;
  signal n_6, n_7, n_8, r1, r2 : std_logic;
  signal r3, r4, r5, r6, r7 : std_logic;
  signal r8, r9, r10 : std_logic;

begin

  g54 : INVD4BWP7T port map(I => vsync, ZN => enable_calc);
  g137 : ND2D4BWP7T port map(A1 => n_8, A2 => n_7, ZN => r);
  g138 : INR3D0BWP7T port map(A1 => n_6, B1 => r3, B2 => r4, ZN => n_8);
  g139 : NR4D0BWP7T port map(A1 => r5, A2 => r6, A3 => r9, A4 => r10, ZN => n_7);
  g140 : NR4D0BWP7T port map(A1 => r7, A2 => r8, A3 => r2, A4 => r1, ZN => n_6);
  g141 : ND2D4BWP7T port map(A1 => n_5, A2 => n_4, ZN => g);
  g142 : INR3D0BWP7T port map(A1 => n_3, B1 => g3, B2 => g4, ZN => n_5);
  g143 : NR4D0BWP7T port map(A1 => g10, A2 => g9, A3 => g6, A4 => g5, ZN => n_4);
  g144 : NR4D0BWP7T port map(A1 => g8, A2 => g7, A3 => g1, A4 => g2, ZN => n_3);
  g145 : ND2D4BWP7T port map(A1 => n_2, A2 => n_1, ZN => b);
  g146 : INR3D0BWP7T port map(A1 => n_0, B1 => b3, B2 => b4, ZN => n_2);
  g147 : NR4D0BWP7T port map(A1 => b10, A2 => b9, A3 => b6, A4 => b5, ZN => n_1);
  g148 : NR4D0BWP7T port map(A1 => b8, A2 => b7, A3 => b2, A4 => b1, ZN => n_0);
  l06_g11912 : OR4D1BWP7T port map(A1 => l06_n_277, A2 => l06_n_295, A3 => l06_n_297, A4 => l06_n_325, Z => g4);
  l06_g11913 : OR2D1BWP7T port map(A1 => l06_n_323, A2 => l06_n_297, Z => r4);
  l06_g11914 : OAI211D1BWP7T port map(A1 => l06_n_114, A2 => l06_n_254, B => l06_n_324, C => l06_n_285, ZN => b4);
  l06_g11915 : OAI211D1BWP7T port map(A1 => l06_n_183, A2 => l06_n_290, B => l06_n_322, C => l06_n_252, ZN => l06_n_325);
  l06_g11916 : AOI31D0BWP7T port map(A1 => l06_n_250, A2 => l06_n_232, A3 => l06_n_160, B => l06_n_321, ZN => l06_n_324);
  l06_g11917 : OAI221D0BWP7T port map(A1 => l06_n_269, A2 => l06_n_122, B1 => l06_n_251, B2 => l06_n_247, C => l06_n_320, ZN => l06_n_323);
  l06_g11918 : NR4D0BWP7T port map(A1 => l06_n_318, A2 => l06_n_304, A3 => l06_n_296, A4 => l06_n_263, ZN => l06_n_322);
  l06_g11919 : OAI211D1BWP7T port map(A1 => l06_n_191, A2 => l06_n_273, B => l06_n_319, C => l06_n_291, ZN => l06_n_321);
  l06_g11920 : NR4D0BWP7T port map(A1 => l06_n_317, A2 => l06_n_304, A3 => l06_n_263, A4 => l06_n_262, ZN => l06_n_320);
  l06_g11921 : NR4D0BWP7T port map(A1 => l06_n_315, A2 => l06_n_275, A3 => l06_n_276, A4 => l06_n_279, ZN => l06_n_319);
  l06_g11922 : OAI221D0BWP7T port map(A1 => l06_n_253, A2 => l06_n_177, B1 => l06_n_202, B2 => l06_n_267, C => l06_n_316, ZN => l06_n_318);
  l06_g11923 : OAI211D1BWP7T port map(A1 => l06_n_162, A2 => l06_n_290, B => l06_n_313, C => l06_n_283, ZN => l06_n_317);
  l06_g11924 : AOI211XD0BWP7T port map(A1 => l06_n_268, A2 => l06_n_198, B => l06_n_312, C => l06_n_262, ZN => l06_n_316);
  l06_g11925 : OAI211D1BWP7T port map(A1 => l06_n_235, A2 => l06_n_251, B => l06_n_314, C => l06_n_299, ZN => l06_n_315);
  l06_g11926 : AOI211XD0BWP7T port map(A1 => l06_n_268, A2 => l06_n_203, B => l06_n_311, C => l06_n_293, ZN => l06_n_314);
  l06_g11927 : AN4D1BWP7T port map(A1 => l06_n_309, A2 => l06_n_306, A3 => l06_n_298, A4 => l06_n_303, Z => l06_n_313);
  l06_g11928 : OAI211D1BWP7T port map(A1 => l06_n_208, A2 => l06_n_280, B => l06_n_308, C => l06_n_300, ZN => l06_n_312);
  l06_g11929 : OAI221D0BWP7T port map(A1 => l06_n_251, A2 => l06_n_241, B1 => l06_n_207, B2 => l06_n_280, C => l06_n_307, ZN => l06_n_311);
  l06_g11930 : IND4D0BWP7T port map(A1 => l06_n_301, B1 => l06_n_254, B2 => l06_n_256, B3 => l06_n_269, ZN => enable4);
  l06_g11931 : NR4D0BWP7T port map(A1 => l06_n_305, A2 => l06_n_296, A3 => l06_n_278, A4 => l06_n_266, ZN => l06_n_309);
  l06_g11932 : AOI222D0BWP7T port map(A1 => l06_n_289, A2 => l06_n_215, B1 => l06_n_288, B2 => l06_n_225, C1 => l06_n_287, C2 => l06_n_210, ZN => l06_n_308);
  l06_g11933 : AOI211XD0BWP7T port map(A1 => l06_n_289, A2 => l06_n_212, B => l06_n_302, C => l06_n_286, ZN => l06_n_307);
  l06_g11934 : AOI21D0BWP7T port map(A1 => l06_n_288, A2 => l06_n_1, B => l06_n_294, ZN => l06_n_306);
  l06_g11935 : IOA21D1BWP7T port map(A1 => l06_n_268, A2 => l06_n_115, B => l06_n_292, ZN => l06_n_305);
  l06_g11936 : AO21D0BWP7T port map(A1 => l06_n_173, A2 => l06_n_177, B => l06_n_280, Z => l06_n_303);
  l06_g11937 : OA31D1BWP7T port map(A1 => l06_n_108, A2 => l06_n_200, A3 => l06_n_214, B => l06_n_287, Z => l06_n_302);
  l06_g11938 : OAI21D0BWP7T port map(A1 => l06_n_265, A2 => l06_n_251, B => l06_n_261, ZN => l06_n_301);
  l06_g11939 : OAI31D0BWP7T port map(A1 => l06_n_83, A2 => l06_n_120, A3 => l06_n_164, B => l06_n_281, ZN => l06_n_300);
  l06_g11940 : IOA21D1BWP7T port map(A1 => l06_n_201, A2 => l06_n_179, B => l06_n_288, ZN => l06_n_299);
  l06_g11941 : OAI21D0BWP7T port map(A1 => l06_n_172, A2 => l06_n_181, B => l06_n_289, ZN => l06_n_298);
  l06_g11942 : OAI211D1BWP7T port map(A1 => l06_n_176, A2 => l06_n_261, B => l06_n_274, C => l06_n_264, ZN => l06_n_304);
  l06_g11943 : OAI22D0BWP7T port map(A1 => l06_n_272, A2 => l06_n_197, B1 => l06_n_269, B2 => l06_n_134, ZN => l06_n_295);
  l06_g11944 : AOI21D0BWP7T port map(A1 => l06_n_183, A2 => l06_n_145, B => l06_n_282, ZN => l06_n_294);
  l06_g11945 : AOI21D0BWP7T port map(A1 => l06_n_184, A2 => l06_n_179, B => l06_n_282, ZN => l06_n_293);
  l06_g11946 : OAI21D0BWP7T port map(A1 => l06_n_195, A2 => l06_n_15, B => l06_n_287, ZN => l06_n_292);
  l06_g11947 : AOI31D0BWP7T port map(A1 => l06_n_250, A2 => l06_n_233, A3 => l06_n_133, B => l06_n_284, ZN => l06_n_291);
  l06_g11948 : NR3D0BWP7T port map(A1 => l06_n_271, A2 => l06_n_59, A3 => l06_n_10, ZN => l06_n_297);
  l06_g11949 : OAI22D0BWP7T port map(A1 => l06_n_253, A2 => l06_n_190, B1 => l06_n_267, B2 => l06_n_2, ZN => l06_n_296);
  l06_g11950 : AOI31D0BWP7T port map(A1 => l06_n_204, A2 => l06_n_199, A3 => l06_n_96, B => l06_n_267, ZN => l06_n_286);
  l06_g11951 : AO21D0BWP7T port map(A1 => l06_n_197, A2 => l06_n_89, B => l06_n_271, Z => l06_n_285);
  l06_g11952 : NR2D0BWP7T port map(A1 => l06_n_269, A2 => l06_n_183, ZN => l06_n_284);
  l06_g11953 : AO21D0BWP7T port map(A1 => l06_n_148, A2 => l06_n_135, B => l06_n_272, Z => l06_n_283);
  l06_g11954 : CKAN2D1BWP7T port map(A1 => l06_n_273, A2 => l06_n_271, Z => l06_n_290);
  l06_g11955 : NR2D1BWP7T port map(A1 => l06_n_270, A2 => l06_n_131, ZN => l06_n_289);
  l06_g11956 : NR2D1BWP7T port map(A1 => l06_n_270, A2 => l06_n_152, ZN => l06_n_288);
  l06_g11957 : NR2D1BWP7T port map(A1 => l06_n_270, A2 => l06_n_150, ZN => l06_n_287);
  l06_g11958 : INVD0BWP7T port map(I => l06_n_282, ZN => l06_n_281);
  l06_g11959 : MOAI22D0BWP7T port map(A1 => l06_n_253, A2 => l06_n_223, B1 => l06_n_257, B2 => l06_n_239, ZN => l06_n_279);
  l06_g11960 : IAO21D0BWP7T port map(A1 => l06_n_194, A2 => l06_n_15, B => l06_n_267, ZN => l06_n_278);
  l06_g11961 : OAI22D0BWP7T port map(A1 => l06_n_258, A2 => l06_n_240, B1 => l06_n_254, B2 => l06_n_84, ZN => l06_n_277);
  l06_g11962 : OAI22D0BWP7T port map(A1 => l06_n_251, A2 => l06_n_246, B1 => l06_n_256, B2 => l06_n_26, ZN => l06_n_276);
  l06_g11963 : AOI21D0BWP7T port map(A1 => l06_n_197, A2 => l06_n_67, B => l06_n_272, ZN => l06_n_275);
  l06_g11964 : AOI32D1BWP7T port map(A1 => l06_n_250, A2 => l06_n_237, A3 => l06_n_78, B1 => l06_n_255, B2 => l06_n_159, ZN => l06_n_274);
  l06_g11965 : ND3D0BWP7T port map(A1 => l06_n_259, A2 => l06_n_140, A3 => l06_n_97, ZN => l06_n_282);
  l06_g11966 : ND3D0BWP7T port map(A1 => l06_n_259, A2 => l06_n_156, A3 => l06_n_97, ZN => l06_n_280);
  l06_g11967 : ND2D1BWP7T port map(A1 => l06_n_260, A2 => l06_n_166, ZN => l06_n_273);
  l06_g11968 : ND2D1BWP7T port map(A1 => l06_n_260, A2 => l06_n_167, ZN => l06_n_272);
  l06_g11969 : ND2D1BWP7T port map(A1 => l06_n_260, A2 => l06_n_147, ZN => l06_n_271);
  l06_g11970 : ND2D1BWP7T port map(A1 => l06_n_259, A2 => l06_n_98, ZN => l06_n_270);
  l06_g11971 : ND2D1BWP7T port map(A1 => l06_n_260, A2 => l06_n_142, ZN => l06_n_269);
  l06_g11972 : IAO21D0BWP7T port map(A1 => l06_n_182, A2 => l06_n_115, B => l06_n_253, ZN => l06_n_266);
  l06_g11973 : NR4D0BWP7T port map(A1 => l06_n_249, A2 => l06_n_237, A3 => l06_n_227, A4 => l06_n_230, ZN => l06_n_265);
  l06_g11974 : OAI211D1BWP7T port map(A1 => l06_n_226, A2 => l06_n_231, B => l06_n_250, C => l06_n_65, ZN => l06_n_264);
  l06_g11975 : AN2D1BWP7T port map(A1 => l06_n_259, A2 => l06_n_174, Z => l06_n_268);
  l06_g11976 : ND3D0BWP7T port map(A1 => l06_n_259, A2 => l06_n_123, A3 => l06_n_372, ZN => l06_n_267);
  l06_g11977 : NR2D1BWP7T port map(A1 => l06_n_251, A2 => l06_n_243, ZN => l06_n_263);
  l06_g11978 : NR3D0BWP7T port map(A1 => l06_n_251, A2 => l06_n_228, A3 => l06_n_189, ZN => l06_n_262);
  l06_g11979 : ND2D1BWP7T port map(A1 => l06_n_250, A2 => l06_n_234, ZN => l06_n_261);
  l06_g11980 : NR2D1BWP7T port map(A1 => l06_n_251, A2 => l06_n_3, ZN => l06_n_260);
  l06_g11981 : NR2D1BWP7T port map(A1 => l06_n_251, A2 => l06_n_221, ZN => l06_n_259);
  l06_g11982 : INVD0BWP7T port map(I => l06_n_257, ZN => l06_n_258);
  l06_g11983 : CKND1BWP7T port map(I => l06_n_255, ZN => l06_n_256);
  l06_g11984 : IND3D1BWP7T port map(A1 => l06_n_114, B1 => l06_n_239, B2 => l06_n_250, ZN => l06_n_252);
  l06_g11985 : AOI21D0BWP7T port map(A1 => l06_n_114, A2 => l06_n_86, B => l06_n_251, ZN => l06_n_257);
  l06_g11986 : NR3D0BWP7T port map(A1 => l06_n_251, A2 => l06_n_220, A3 => l06_n_149, ZN => l06_n_255);
  l06_g11987 : ND4D0BWP7T port map(A1 => l06_n_250, A2 => l06_n_213, A3 => l06_n_174, A4 => l06_n_101, ZN => l06_n_254);
  l06_g11988 : ND3D0BWP7T port map(A1 => l06_n_250, A2 => l06_n_209, A3 => l06_n_42, ZN => l06_n_253);
  l06_g11989 : INVD1BWP7T port map(I => l06_n_251, ZN => l06_n_250);
  l06_g11990 : OAI211D1BWP7T port map(A1 => l06_n_25, A2 => l06_n_53, B => l06_n_248, C => l06_n_109, ZN => l06_n_251);
  l06_g11991 : ND3D0BWP7T port map(A1 => l06_n_245, A2 => l06_n_242, A3 => l06_n_221, ZN => l06_n_249);
  l06_g11992 : AOI211D1BWP7T port map(A1 => l06_n_38, A2 => l06_n_37, B => l06_n_244, C => l06_n_236, ZN => l06_n_248);
  l06_g11993 : OA22D0BWP7T port map(A1 => l06_n_245, A2 => l06_n_77, B1 => l06_n_86, B2 => l06_n_240, Z => l06_n_247);
  l06_g11994 : AOI222D0BWP7T port map(A1 => l06_n_227, A2 => l06_n_187, B1 => l06_n_230, B2 => l06_n_185, C1 => l06_n_226, C2 => l06_n_161, ZN => l06_n_246);
  l06_g11995 : OAI22D0BWP7T port map(A1 => l06_n_229, A2 => l06_n_168, B1 => l06_n_38, B2 => l06_n_37, ZN => l06_n_244);
  l06_g11996 : INR2D1BWP7T port map(A1 => l06_n_240, B1 => l06_n_239, ZN => l06_n_245);
  l06_g11997 : AOI22D0BWP7T port map(A1 => l06_n_230, A2 => l06_n_139, B1 => l06_n_227, B2 => l06_n_111, ZN => l06_n_243);
  l06_g11998 : NR3D0BWP7T port map(A1 => l06_n_226, A2 => l06_n_231, A3 => l06_n_224, ZN => l06_n_242);
  l06_g11999 : AOI21D0BWP7T port map(A1 => l06_n_234, A2 => l06_n_180, B => l06_n_238, ZN => l06_n_241);
  l06_g12000 : IAO21D0BWP7T port map(A1 => l06_n_180, A2 => l06_n_88, B => l06_n_228, ZN => l06_n_238);
  l06_g12001 : NR2XD0BWP7T port map(A1 => l06_n_232, A2 => l06_n_233, ZN => l06_n_240);
  l06_g12002 : OAI22D0BWP7T port map(A1 => l06_n_3, A2 => l06_n_175, B1 => l06_n_217, B2 => l06_n_41, ZN => l06_n_239);
  l06_g12003 : MOAI22D0BWP7T port map(A1 => x(8), A2 => l06_n_9, B1 => l06_n_218, B2 => l06_n_168, ZN => l06_n_236);
  l06_g12004 : AOI31D0BWP7T port map(A1 => l06_n_219, A2 => l06_n_193, A3 => l06_n_141, B => l06_n_222, ZN => l06_n_235);
  l06_g12005 : IOA21D1BWP7T port map(A1 => l06_n_219, A2 => l06_n_167, B => l06_n_5, ZN => l06_n_237);
  l06_g12006 : NR2D1BWP7T port map(A1 => l06_n_216, A2 => l06_n_151, ZN => l06_n_229);
  l06_g12007 : NR2D1BWP7T port map(A1 => l06_n_220, A2 => l06_n_175, ZN => l06_n_234);
  l06_g12008 : NR2XD0BWP7T port map(A1 => l06_n_3, A2 => l06_n_149, ZN => l06_n_233);
  l06_g12009 : NR2XD0BWP7T port map(A1 => l06_n_3, A2 => l06_n_171, ZN => l06_n_232);
  l06_g12010 : INR2D1BWP7T port map(A1 => l06_n_147, B1 => l06_n_220, ZN => l06_n_231);
  l06_g12011 : NR2D1BWP7T port map(A1 => l06_n_220, A2 => l06_n_171, ZN => l06_n_230);
  l06_g12012 : ND4D0BWP7T port map(A1 => l06_n_204, A2 => l06_n_75, A3 => l06_n_77, A4 => l06_n_13, ZN => l06_n_225);
  l06_g12013 : IAO21D0BWP7T port map(A1 => l06_n_193, A2 => l06_n_166, B => l06_n_3, ZN => l06_n_224);
  l06_g12014 : NR3D0BWP7T port map(A1 => l06_n_214, A2 => l06_n_157, A3 => l06_n_146, ZN => l06_n_223);
  l06_g12015 : IAO21D0BWP7T port map(A1 => l06_n_90, A2 => l06_n_65, B => l06_n_5, ZN => l06_n_222);
  l06_g12016 : IND4D0BWP7T port map(A1 => l06_n_41, B1 => l06_n_99, B2 => l06_n_107, B3 => l06_n_211, ZN => l06_n_228);
  l06_g12017 : INR2D1BWP7T port map(A1 => l06_n_142, B1 => l06_n_220, ZN => l06_n_227);
  l06_g12018 : INR2D1BWP7T port map(A1 => l06_n_166, B1 => l06_n_220, ZN => l06_n_226);
  l06_g12019 : INVD0BWP7T port map(I => l06_n_220, ZN => l06_n_219);
  l06_g12020 : OAI222D0BWP7T port map(A1 => l06_n_205, A2 => l06_n_151, B1 => l06_n_29, B2 => l06_n_49, C1 => l06_n_92, C2 => l06_n_47, ZN => l06_n_218);
  l06_g12021 : IND2D1BWP7T port map(A1 => l06_n_101, B1 => l06_n_211, ZN => l06_n_221);
  l06_g12023 : ND2D1BWP7T port map(A1 => l06_n_211, A2 => l06_n_100, ZN => l06_n_220);
  l06_g12024 : IND3D1BWP7T port map(A1 => l06_n_107, B1 => l06_n_99, B2 => l06_n_213, ZN => l06_n_217);
  l06_g12025 : OAI222D0BWP7T port map(A1 => l06_n_196, A2 => l06_n_116, B1 => x(5), B2 => l06_n_112, C1 => l06_n_28, C2 => l06_n_47, ZN => l06_n_216);
  l06_g12026 : ND4D0BWP7T port map(A1 => l06_n_201, A2 => l06_n_155, A3 => l06_n_76, A4 => l06_n_64, ZN => l06_n_215);
  l06_g12029 : IND2D1BWP7T port map(A1 => l06_n_181, B1 => l06_n_207, ZN => l06_n_212);
  l06_g12030 : ND2D1BWP7T port map(A1 => l06_n_204, A2 => l06_n_70, ZN => l06_n_214);
  l06_g12031 : AOI211D1BWP7T port map(A1 => l06_n_43, A2 => l06_n_23, B => l06_n_206, C => l06_n_72, ZN => l06_n_213);
  l06_g12032 : OR3D1BWP7T port map(A1 => l06_n_128, A2 => l06_n_188, A3 => l06_n_195, Z => l06_n_210);
  l06_g12033 : AOI211D1BWP7T port map(A1 => l06_n_154, A2 => y(4), B => l06_n_163, C => l06_n_206, ZN => l06_n_209);
  l06_g12034 : INR4D0BWP7T port map(A1 => l06_n_155, B1 => l06_n_60, B2 => l06_n_158, B3 => l06_n_194, ZN => l06_n_208);
  l06_g12035 : AOI211D1BWP7T port map(A1 => l06_n_43, A2 => l06_n_31, B => l06_n_206, C => l06_n_73, ZN => l06_n_211);
  l06_g12036 : OAI21D0BWP7T port map(A1 => l06_n_170, A2 => l06_n_116, B => l06_n_117, ZN => l06_n_205);
  l06_g12037 : AN3D1BWP7T port map(A1 => l06_n_186, A2 => l06_n_184, A3 => l06_n_135, Z => l06_n_207);
  l06_g12038 : ND3D0BWP7T port map(A1 => l06_n_169, A2 => l06_n_143, A3 => l06_n_130, ZN => l06_n_206);
  l06_g12039 : AO21D0BWP7T port map(A1 => l06_n_85, A2 => l06_n_11, B => l06_n_198, Z => l06_n_203);
  l06_g12040 : AOI211XD0BWP7T port map(A1 => l06_n_118, A2 => l06_n_12, B => l06_n_188, C => l06_n_178, ZN => l06_n_202);
  l06_g12041 : INR3D0BWP7T port map(A1 => l06_n_67, B1 => l06_n_44, B2 => l06_n_182, ZN => l06_n_204);
  l06_g12042 : INVD0BWP7T port map(I => l06_n_199, ZN => l06_n_200);
  l06_g12043 : AN2D0BWP7T port map(A1 => l06_n_170, A2 => l06_n_117, Z => l06_n_196);
  l06_g12044 : INR2XD0BWP7T port map(A1 => l06_n_184, B1 => l06_n_181, ZN => l06_n_201);
  l06_g12045 : NR2XD0BWP7T port map(A1 => l06_n_185, A2 => l06_n_71, ZN => l06_n_199);
  l06_g12046 : ND2D1BWP7T port map(A1 => l06_n_189, A2 => l06_n_76, ZN => l06_n_198);
  l06_g12047 : NR2XD0BWP7T port map(A1 => l06_n_178, A2 => l06_n_44, ZN => l06_n_197);
  l06_g12048 : OA21D0BWP7T port map(A1 => l06_n_46, A2 => l06_n_6, B => l06_n_169, Z => l06_n_192);
  l06_g12049 : AOI21D0BWP7T port map(A1 => l06_n_66, A2 => l06_n_11, B => l06_n_178, ZN => l06_n_191);
  l06_g12050 : INR3D0BWP7T port map(A1 => l06_n_89, B1 => l06_n_44, B2 => l06_n_157, ZN => l06_n_190);
  l06_g12051 : ND4D0BWP7T port map(A1 => l06_n_2, A2 => l06_n_74, A3 => l06_n_84, A4 => l06_n_67, ZN => l06_n_195);
  l06_g12052 : IND2D1BWP7T port map(A1 => l06_n_182, B1 => l06_n_114, ZN => l06_n_194);
  l06_g12053 : OR2D1BWP7T port map(A1 => l06_n_167, A2 => l06_n_147, Z => l06_n_193);
  l06_g12054 : INVD0BWP7T port map(I => l06_n_186, ZN => l06_n_187);
  l06_g12055 : INVD0BWP7T port map(I => l06_n_180, ZN => l06_n_179);
  l06_g12056 : CKND1BWP7T port map(I => l06_n_178, ZN => l06_n_177);
  l06_g12057 : INR2XD0BWP7T port map(A1 => l06_n_86, B1 => l06_n_146, ZN => l06_n_176);
  l06_g12058 : NR2XD0BWP7T port map(A1 => l06_n_146, A2 => l06_n_61, ZN => l06_n_189);
  l06_g12059 : IND2D1BWP7T port map(A1 => l06_n_71, B1 => l06_n_145, ZN => l06_n_188);
  l06_g12060 : NR2XD0BWP7T port map(A1 => l06_n_161, A2 => l06_n_83, ZN => l06_n_186);
  l06_g12061 : OR2D1BWP7T port map(A1 => l06_n_146, A2 => l06_n_65, Z => l06_n_185);
  l06_g12062 : CKAN2D1BWP7T port map(A1 => l06_n_148, A2 => l06_n_89, Z => l06_n_184);
  l06_g12063 : NR2XD0BWP7T port map(A1 => l06_n_160, A2 => l06_n_88, ZN => l06_n_183);
  l06_g12064 : ND2D1BWP7T port map(A1 => l06_n_153, A2 => l06_n_62, ZN => l06_n_182);
  l06_g12065 : OR2D1BWP7T port map(A1 => l06_n_158, A2 => l06_n_12, Z => l06_n_181);
  l06_g12066 : IND2D1BWP7T port map(A1 => l06_n_159, B1 => l06_n_135, ZN => l06_n_180);
  l06_g12067 : ND2D1BWP7T port map(A1 => l06_n_153, A2 => l06_n_134, ZN => l06_n_178);
  l06_g12068 : CKND1BWP7T port map(I => l06_n_172, ZN => l06_n_173);
  l06_g12069 : NR4D0BWP7T port map(A1 => l06_n_128, A2 => l06_n_120, A3 => l06_n_108, A4 => l06_n_82, ZN => l06_n_165);
  l06_g12070 : OAI211D1BWP7T port map(A1 => l06_n_13, A2 => l06_n_59, B => l06_n_162, C => l06_n_91, ZN => l06_n_164);
  l06_g12071 : IAO21D0BWP7T port map(A1 => l06_n_136, A2 => l06_n_43, B => y(4), ZN => l06_n_163);
  l06_g12072 : OR2D1BWP7T port map(A1 => l06_n_152, A2 => l06_n_98, Z => l06_n_175);
  l06_g12073 : INR2D1BWP7T port map(A1 => l06_n_97, B1 => l06_n_4, ZN => l06_n_174);
  l06_g12074 : OAI211D1BWP7T port map(A1 => l06_n_14, A2 => l06_n_68, B => l06_n_145, C => l06_n_138, ZN => l06_n_172);
  l06_g12075 : OR2D1BWP7T port map(A1 => l06_n_150, A2 => l06_n_98, Z => l06_n_171);
  l06_g12076 : AO21D0BWP7T port map(A1 => l06_n_50, A2 => x(2), B => l06_n_144, Z => l06_n_170);
  l06_g12077 : AOI211XD0BWP7T port map(A1 => l06_n_35, A2 => y(9), B => l06_n_124, C => l06_n_127, ZN => l06_n_169);
  l06_g12078 : OAI22D0BWP7T port map(A1 => l06_n_126, A2 => l06_n_49, B1 => l06_n_92, B2 => l06_n_29, ZN => l06_n_168);
  l06_g12079 : NR2D1BWP7T port map(A1 => l06_n_4, A2 => l06_n_97, ZN => l06_n_167);
  l06_g12080 : INR2D1BWP7T port map(A1 => l06_n_156, B1 => l06_n_97, ZN => l06_n_166);
  l06_g12082 : INR2XD0BWP7T port map(A1 => l06_n_135, B1 => l06_n_88, ZN => l06_n_162);
  l06_g12083 : IND2D1BWP7T port map(A1 => l06_n_141, B1 => l06_n_75, ZN => l06_n_161);
  l06_g12084 : ND2D1BWP7T port map(A1 => l06_n_134, A2 => l06_n_76, ZN => l06_n_160);
  l06_g12085 : OR2D1BWP7T port map(A1 => l06_n_139, A2 => l06_n_83, Z => l06_n_159);
  l06_g12086 : OAI21D0BWP7T port map(A1 => l06_n_110, A2 => l06_n_13, B => l06_n_91, ZN => l06_n_158);
  l06_g12087 : IND2D1BWP7T port map(A1 => l06_n_128, B1 => l06_n_93, ZN => l06_n_157);
  l06_g12088 : NR2D1BWP7T port map(A1 => l06_n_129, A2 => l06_n_104, ZN => l06_n_156);
  l06_g12089 : CKAN2D1BWP7T port map(A1 => l06_n_132, A2 => l06_n_138, Z => l06_n_155);
  l06_g12090 : IND2D1BWP7T port map(A1 => l06_n_136, B1 => l06_n_43, ZN => l06_n_154);
  l06_g12091 : INR2XD0BWP7T port map(A1 => l06_n_76, B1 => l06_n_125, ZN => l06_n_153);
  l06_g12092 : MAOI222D1BWP7T port map(A => l06_n_95, B => x(2), C => x_player(2), ZN => l06_n_144);
  l06_g12093 : AOI22D0BWP7T port map(A1 => l06_n_113, A2 => y(5), B1 => l06_n_46, B2 => y_player(5), ZN => l06_n_143);
  l06_g12094 : IND2D1BWP7T port map(A1 => l06_n_129, B1 => l06_n_104, ZN => l06_n_152);
  l06_g12096 : NR3D0BWP7T port map(A1 => l06_n_116, A2 => l06_n_50, A3 => x(2), ZN => l06_n_151);
  l06_g12097 : ND2D1BWP7T port map(A1 => l06_n_137, A2 => l06_n_105, ZN => l06_n_150);
  l06_g12098 : OR2D1BWP7T port map(A1 => l06_n_131, A2 => l06_n_98, Z => l06_n_149);
  l06_g12099 : OAI21D0BWP7T port map(A1 => l06_n_118, A2 => l06_n_57, B => l06_n_11, ZN => l06_n_148);
  l06_g12100 : INR2D1BWP7T port map(A1 => l06_n_140, B1 => l06_n_97, ZN => l06_n_147);
  l06_g12101 : ND3D0BWP7T port map(A1 => l06_n_114, A2 => l06_n_75, A3 => l06_n_79, ZN => l06_n_146);
  l06_g12102 : OA21D0BWP7T port map(A1 => l06_n_59, A2 => l06_n_14, B => l06_n_132, Z => l06_n_145);
  l06_g12103 : INVD1BWP7T port map(I => l06_n_133, ZN => l06_n_134);
  l06_g12104 : INR2D1BWP7T port map(A1 => l06_n_123, B1 => l06_n_372, ZN => l06_n_142);
  l06_g12105 : ND2D1BWP7T port map(A1 => l06_n_119, A2 => l06_n_121, ZN => l06_n_141);
  l06_g12106 : NR2D1BWP7T port map(A1 => l06_n_371, A2 => l06_n_80, ZN => l06_n_140);
  l06_g12107 : ND2D1BWP7T port map(A1 => l06_n_121, A2 => l06_n_75, ZN => l06_n_139);
  l06_g12108 : CKAN2D1BWP7T port map(A1 => l06_n_119, A2 => l06_n_75, Z => l06_n_138);
  l06_g12109 : NR2D1BWP7T port map(A1 => l06_n_106, A2 => l06_n_48, ZN => l06_n_137);
  l06_g12110 : ND2D1BWP7T port map(A1 => l06_n_99, A2 => l06_n_41, ZN => l06_n_136);
  l06_g12111 : CKAN2D1BWP7T port map(A1 => l06_n_122, A2 => l06_n_76, Z => l06_n_135);
  l06_g12112 : ND2D1BWP7T port map(A1 => l06_n_114, A2 => l06_n_62, ZN => l06_n_133);
  l06_g12113 : MOAI22D0BWP7T port map(A1 => l06_n_35, A2 => y(9), B1 => l06_n_46, B2 => l06_n_6, ZN => l06_n_127);
  l06_g12114 : AN3D0BWP7T port map(A1 => l06_n_47, A2 => l06_n_92, A3 => l06_n_29, Z => l06_n_126);
  l06_g12115 : OA21D0BWP7T port map(A1 => l06_n_85, A2 => l06_n_60, B => l06_n_11, Z => l06_n_125);
  l06_g12116 : MOAI22D0BWP7T port map(A1 => l06_n_52, A2 => l06_n_24, B1 => l06_n_52, B2 => l06_n_24, ZN => l06_n_124);
  l06_g12118 : AOI21D0BWP7T port map(A1 => l06_n_57, A2 => l06_n_15, B => l06_n_115, ZN => l06_n_132);
  l06_g12119 : IND2D1BWP7T port map(A1 => l06_n_80, B1 => l06_n_371, ZN => l06_n_131);
  l06_g12120 : MOAI22D0BWP7T port map(A1 => l06_n_54, A2 => l06_n_34, B1 => l06_n_54, B2 => l06_n_34, ZN => l06_n_130);
  l06_g12121 : IND2D1BWP7T port map(A1 => l06_n_48, B1 => l06_n_106, ZN => l06_n_129);
  l06_g12122 : AOI21D0BWP7T port map(A1 => l06_n_87, A2 => l06_n_59, B => l06_n_13, ZN => l06_n_128);
  l06_g12123 : NR2D1BWP7T port map(A1 => l06_n_46, A2 => y_player(5), ZN => l06_n_113);
  l06_g12124 : ND2D1BWP7T port map(A1 => l06_n_49, A2 => x_player(5), ZN => l06_n_112);
  l06_g12125 : IND2D1BWP7T port map(A1 => l06_n_65, B1 => l06_n_79, ZN => l06_n_111);
  l06_g12126 : NR2XD0BWP7T port map(A1 => l06_n_85, A2 => l06_n_63, ZN => l06_n_110);
  l06_g12127 : ND2D1BWP7T port map(A1 => l06_n_53, A2 => l06_n_25, ZN => l06_n_109);
  l06_g12128 : NR2D1BWP7T port map(A1 => l06_n_81, A2 => l06_n_56, ZN => l06_n_123);
  l06_g12129 : CKAN2D1BWP7T port map(A1 => l06_n_77, A2 => l06_n_62, Z => l06_n_122);
  l06_g12130 : ND2D1BWP7T port map(A1 => l06_n_85, A2 => l06_n_27, ZN => l06_n_121);
  l06_g12131 : ND2D1BWP7T port map(A1 => l06_n_75, A2 => l06_n_70, ZN => l06_n_120);
  l06_g12132 : NR2XD0BWP7T port map(A1 => l06_n_78, A2 => l06_n_90, ZN => l06_n_119);
  l06_g12133 : IND2D1BWP7T port map(A1 => l06_n_85, B1 => l06_n_87, ZN => l06_n_118);
  l06_g12134 : ND2D1BWP7T port map(A1 => l06_n_51, A2 => l06_n_33, ZN => l06_n_117);
  l06_g12135 : NR2XD0BWP7T port map(A1 => l06_n_51, A2 => l06_n_33, ZN => l06_n_116);
  l06_g12136 : NR2D1BWP7T port map(A1 => l06_n_87, A2 => l06_n_14, ZN => l06_n_115);
  l06_g12137 : CKAN2D1BWP7T port map(A1 => l06_n_84, A2 => l06_n_77, Z => l06_n_114);
  l06_g12140 : OAI21D0BWP7T port map(A1 => l06_n_57, A2 => l06_n_63, B => l06_n_12, ZN => l06_n_96);
  l06_g12141 : AOI22D0BWP7T port map(A1 => l06_n_39, A2 => x(0), B1 => x(1), B2 => l06_n_7, ZN => l06_n_95);
  l06_g12143 : OAI21D0BWP7T port map(A1 => l06_n_57, A2 => l06_n_69, B => l06_n_12, ZN => l06_n_93);
  l06_g12144 : AOI21D0BWP7T port map(A1 => l06_n_0, A2 => l06_n_16, B => l06_n_13, ZN => l06_n_108);
  l06_g12145 : MAOI22D0BWP7T port map(A1 => l06_n_42, A2 => y(3), B1 => l06_n_42, B2 => y(3), ZN => l06_n_107);
  l06_g12146 : MOAI22D0BWP7T port map(A1 => l06_n_45, A2 => y(0), B1 => l06_n_45, B2 => y(0), ZN => l06_n_106);
  l06_g12147 : MOAI22D0BWP7T port map(A1 => l06_n_56, A2 => l06_n_18, B1 => l06_n_56, B2 => l06_n_18, ZN => l06_n_105);
  l06_g12148 : MAOI22D0BWP7T port map(A1 => l06_n_56, A2 => l06_n_30, B1 => l06_n_56, B2 => l06_n_30, ZN => l06_n_104);
  l06_g12151 : MOAI22D0BWP7T port map(A1 => l06_n_42, A2 => l06_n_32, B1 => l06_n_42, B2 => l06_n_32, ZN => l06_n_101);
  l06_g12152 : MAOI22D0BWP7T port map(A1 => l06_n_42, A2 => l06_n_21, B1 => l06_n_42, B2 => l06_n_21, ZN => l06_n_100);
  l06_g12153 : INR2D1BWP7T port map(A1 => l06_n_56, B1 => l06_n_81, ZN => l06_n_99);
  l06_g12154 : MAOI22D0BWP7T port map(A1 => l06_n_41, A2 => l06_n_20, B1 => l06_n_41, B2 => l06_n_20, ZN => l06_n_98);
  l06_g12155 : MAOI22D0BWP7T port map(A1 => l06_n_41, A2 => l06_n_22, B1 => l06_n_41, B2 => l06_n_22, ZN => l06_n_97);
  l06_g12156 : INVD1BWP7T port map(I => l06_n_28, ZN => l06_n_92);
  l06_g12157 : INVD0BWP7T port map(I => l06_n_84, ZN => l06_n_83);
  l06_g12158 : NR2D0BWP7T port map(A1 => l06_n_64, A2 => l06_n_26, ZN => l06_n_82);
  l06_g12159 : OR2D1BWP7T port map(A1 => l06_n_64, A2 => l06_n_10, Z => l06_n_91);
  l06_g12160 : NR2D0BWP7T port map(A1 => l06_n_64, A2 => l06_n_14, ZN => l06_n_90);
  l06_g12161 : ND2D1BWP7T port map(A1 => l06_n_69, A2 => l06_n_11, ZN => l06_n_89);
  l06_g12162 : NR2D0BWP7T port map(A1 => l06_n_68, A2 => l06_n_10, ZN => l06_n_88);
  l06_g12163 : NR2XD0BWP7T port map(A1 => l06_n_60, A2 => l06_n_66, ZN => l06_n_87);
  l06_g12164 : ND2D1BWP7T port map(A1 => l06_n_69, A2 => l06_n_27, ZN => l06_n_86);
  l06_g12165 : ND2D1BWP7T port map(A1 => l06_n_59, A2 => l06_n_68, ZN => l06_n_85);
  l06_g12166 : ND2D1BWP7T port map(A1 => l06_n_66, A2 => l06_n_27, ZN => l06_n_84);
  l06_g12168 : CKND2D0BWP7T port map(A1 => l06_n_60, A2 => l06_n_11, ZN => l06_n_74);
  l06_g12169 : NR2XD0BWP7T port map(A1 => l06_n_43, A2 => l06_n_31, ZN => l06_n_73);
  l06_g12170 : NR2D1BWP7T port map(A1 => l06_n_43, A2 => l06_n_23, ZN => l06_n_72);
  l06_g12171 : IND2D1BWP7T port map(A1 => l06_n_45, B1 => l06_n_48, ZN => l06_n_81);
  l06_g12172 : CKND2D1BWP7T port map(A1 => l06_n_48, A2 => l06_n_45, ZN => l06_n_80);
  l06_g12173 : ND2D1BWP7T port map(A1 => l06_n_58, A2 => l06_n_27, ZN => l06_n_79);
  l06_g12174 : AN2D1BWP7T port map(A1 => l06_n_63, A2 => l06_n_27, Z => l06_n_78);
  l06_g12175 : ND2D1BWP7T port map(A1 => l06_n_57, A2 => l06_n_27, ZN => l06_n_77);
  l06_g12176 : ND2D1BWP7T port map(A1 => l06_n_63, A2 => l06_n_11, ZN => l06_n_76);
  l06_g12177 : ND2D1BWP7T port map(A1 => l06_n_60, A2 => l06_n_27, ZN => l06_n_75);
  l06_g12178 : INVD1BWP7T port map(I => l06_n_61, ZN => l06_n_62);
  l06_g12179 : INVD1BWP7T port map(I => l06_n_58, ZN => l06_n_59);
  l06_g12180 : INVD1BWP7T port map(I => l06_n_0, ZN => l06_n_57);
  l06_g12182 : NR2D0BWP7T port map(A1 => l06_n_14, A2 => l06_n_16, ZN => l06_n_71);
  l06_g12183 : CKND2D1BWP7T port map(A1 => l06_n_17, A2 => l06_n_12, ZN => l06_n_70);
  l06_g12184 : NR2D0BWP7T port map(A1 => l06_n_16, A2 => draw_count4(0), ZN => l06_n_69);
  l06_g12185 : ND2D1BWP7T port map(A1 => l06_n_17, A2 => draw_count4(0), ZN => l06_n_68);
  l06_g12186 : IND2D1BWP7T port map(A1 => l06_n_16, B1 => l06_n_11, ZN => l06_n_67);
  l06_g12187 : NR2D0BWP7T port map(A1 => l06_n_19, A2 => draw_count4(0), ZN => l06_n_66);
  l06_g12188 : INR2D1BWP7T port map(A1 => l06_n_17, B1 => l06_n_26, ZN => l06_n_65);
  l06_g12189 : IND2D1BWP7T port map(A1 => l06_n_16, B1 => draw_count4(0), ZN => l06_n_64);
  l06_g12190 : INR2D1BWP7T port map(A1 => l06_n_17, B1 => draw_count4(0), ZN => l06_n_63);
  l06_g12191 : NR2D0BWP7T port map(A1 => l06_n_26, A2 => l06_n_16, ZN => l06_n_61);
  l06_g12192 : INR2D1BWP7T port map(A1 => draw_count4(0), B1 => l06_n_36, ZN => l06_n_60);
  l06_g12193 : NR2D0BWP7T port map(A1 => l06_n_36, A2 => draw_count4(0), ZN => l06_n_58);
  l06_g12195 : INR2XD0BWP7T port map(A1 => l06_n_22, B1 => l06_n_20, ZN => l06_n_56);
  l06_g12198 : IAO21D0BWP7T port map(A1 => x(1), A2 => l06_n_7, B => x_player(0), ZN => l06_n_39);
  l06_g12199 : MOAI22D0BWP7T port map(A1 => y(7), A2 => y_player(7), B1 => y(7), B2 => y_player(7), ZN => l06_n_54);
  l06_g12200 : MOAI22D0BWP7T port map(A1 => x(7), A2 => x_player(7), B1 => x(7), B2 => x_player(7), ZN => l06_n_53);
  l06_g12201 : MOAI22D0BWP7T port map(A1 => y(8), A2 => y_player(8), B1 => y(8), B2 => y_player(8), ZN => l06_n_52);
  l06_g12202 : OA21D0BWP7T port map(A1 => l06_n_8, A2 => x_player(4), B => l06_n_28, Z => l06_n_51);
  l06_g12203 : MAOI22D0BWP7T port map(A1 => x(3), A2 => x_player(3), B1 => x(3), B2 => x_player(3), ZN => l06_n_50);
  l06_g12204 : MAOI22D0BWP7T port map(A1 => x(6), A2 => x_player(6), B1 => x(6), B2 => x_player(6), ZN => l06_n_49);
  l06_g12205 : XNR2D1BWP7T port map(A1 => y(0), A2 => y_player(0), ZN => l06_n_48);
  l06_g12206 : MAOI22D0BWP7T port map(A1 => x(5), A2 => x_player(5), B1 => x(5), B2 => x_player(5), ZN => l06_n_47);
  l06_g12207 : MOAI22D0BWP7T port map(A1 => y(6), A2 => y_player(6), B1 => y(6), B2 => y_player(6), ZN => l06_n_46);
  l06_g12208 : OR2D1BWP7T port map(A1 => l06_n_18, A2 => l06_n_30, Z => l06_n_45);
  l06_g12209 : NR2D1BWP7T port map(A1 => l06_n_10, A2 => l06_n_19, ZN => l06_n_44);
  l06_g12210 : MAOI22D0BWP7T port map(A1 => y(5), A2 => y_player(5), B1 => y(5), B2 => y_player(5), ZN => l06_n_43);
  l06_g12211 : IND2D1BWP7T port map(A1 => l06_n_31, B1 => l06_n_23, ZN => l06_n_42);
  l06_g12212 : INR2XD0BWP7T port map(A1 => l06_n_21, B1 => l06_n_32, ZN => l06_n_41);
  l06_g12213 : INVD1BWP7T port map(I => l06_n_27, ZN => l06_n_26);
  l06_g12214 : AN2D1BWP7T port map(A1 => x(8), A2 => l06_n_9, Z => l06_n_38);
  l06_g12215 : IND2D1BWP7T port map(A1 => x(7), B1 => x_player(7), ZN => l06_n_37);
  l06_g12216 : IND2D1BWP7T port map(A1 => draw_count4(2), B1 => draw_count4(1), ZN => l06_n_36);
  l06_g12217 : IND2D1BWP7T port map(A1 => y(8), B1 => y_player(8), ZN => l06_n_35);
  l06_g12218 : IND2D1BWP7T port map(A1 => y(6), B1 => y_player(6), ZN => l06_n_34);
  l06_g12219 : INR2XD0BWP7T port map(A1 => x_player(3), B1 => x(3), ZN => l06_n_33);
  l06_g12220 : INR2D1BWP7T port map(A1 => y(3), B1 => y_player(3), ZN => l06_n_32);
  l06_g12221 : INR2XD0BWP7T port map(A1 => y_player(4), B1 => y(4), ZN => l06_n_31);
  l06_g12222 : INR2XD0BWP7T port map(A1 => y(1), B1 => y_player(1), ZN => l06_n_30);
  l06_g12223 : IND2D1BWP7T port map(A1 => x_player(5), B1 => x(5), ZN => l06_n_29);
  l06_g12224 : ND2D1BWP7T port map(A1 => l06_n_8, A2 => x_player(4), ZN => l06_n_28);
  l06_g12225 : INR2D1BWP7T port map(A1 => draw_count4(3), B1 => draw_count4(4), ZN => l06_n_27);
  l06_g12227 : INVD1BWP7T port map(I => l06_n_15, ZN => l06_n_14);
  l06_g12228 : INVD1BWP7T port map(I => l06_n_13, ZN => l06_n_12);
  l06_g12229 : INVD1BWP7T port map(I => l06_n_11, ZN => l06_n_10);
  l06_g12230 : IND2D1BWP7T port map(A1 => x_player(6), B1 => x(6), ZN => l06_n_25);
  l06_g12231 : INR2D1BWP7T port map(A1 => y_player(7), B1 => y(7), ZN => l06_n_24);
  l06_g12232 : IND2D1BWP7T port map(A1 => y_player(4), B1 => y(4), ZN => l06_n_23);
  l06_g12233 : IND2D1BWP7T port map(A1 => y(2), B1 => y_player(2), ZN => l06_n_22);
  l06_g12234 : IND2D1BWP7T port map(A1 => y(3), B1 => y_player(3), ZN => l06_n_21);
  l06_g12235 : INR2D1BWP7T port map(A1 => y(2), B1 => y_player(2), ZN => l06_n_20);
  l06_g12236 : IND2D1BWP7T port map(A1 => draw_count4(1), B1 => draw_count4(2), ZN => l06_n_19);
  l06_g12237 : INR2XD0BWP7T port map(A1 => y_player(1), B1 => y(1), ZN => l06_n_18);
  l06_g12238 : NR2D0BWP7T port map(A1 => draw_count4(2), A2 => draw_count4(1), ZN => l06_n_17);
  l06_g12239 : ND2D1BWP7T port map(A1 => draw_count4(2), A2 => draw_count4(1), ZN => l06_n_16);
  l06_g12240 : NR2D0BWP7T port map(A1 => draw_count4(4), A2 => draw_count4(3), ZN => l06_n_15);
  l06_g12241 : CKND2D1BWP7T port map(A1 => draw_count4(4), A2 => draw_count4(3), ZN => l06_n_13);
  l06_g12242 : INR2D1BWP7T port map(A1 => draw_count4(4), B1 => draw_count4(3), ZN => l06_n_11);
  l06_g12243 : INVD0BWP7T port map(I => x_player(8), ZN => l06_n_9);
  l06_g12244 : CKND1BWP7T port map(I => x(4), ZN => l06_n_8);
  l06_g12245 : INVD0BWP7T port map(I => x_player(1), ZN => l06_n_7);
  l06_g12246 : INVD1BWP7T port map(I => y(5), ZN => l06_n_6);
  l06_g2 : IIND4D0BWP7T port map(A1 => l06_n_154, A2 => l06_n_42, B1 => l06_n_130, B2 => l06_n_192, ZN => l06_n_5);
  l06_g12247 : IND2D1BWP7T port map(A1 => l06_n_105, B1 => l06_n_137, ZN => l06_n_4);
  l06_g12248 : IND2D1BWP7T port map(A1 => l06_n_100, B1 => l06_n_213, ZN => l06_n_3);
  l06_g12249 : INR3D0BWP7T port map(A1 => l06_n_75, B1 => l06_n_78, B2 => l06_n_44, ZN => l06_n_2);
  l06_g12250 : IND4D0BWP7T port map(A1 => l06_n_44, B1 => l06_n_165, B2 => l06_n_145, B3 => l06_n_153, ZN => l06_n_1);
  l06_g12251 : IND2D1BWP7T port map(A1 => l06_n_19, B1 => draw_count4(0), ZN => l06_n_0);
  l06_g12253 : CKXOR2D1BWP7T port map(A1 => l06_n_56, A2 => y(1), Z => l06_n_371);
  l06_g12254 : CKXOR2D1BWP7T port map(A1 => l06_n_41, A2 => y(2), Z => l06_n_372);
  l042_count_reg_2 : DFCNQD1BWP7T port map(CDN => l042_n_0, CP => clk, D => l042_n_6, Q => draw_count2(2));
  l042_g59 : CKAN2D1BWP7T port map(A1 => enable2, A2 => l042_n_5, Z => l042_n_6);
  l042_count_reg_1 : DFCNQD1BWP7T port map(CDN => l042_n_0, CP => clk, D => l042_n_4, Q => draw_count2(1));
  l042_g61 : MOAI22D0BWP7T port map(A1 => l042_n_1, A2 => draw_count2(2), B1 => l042_n_1, B2 => draw_count2(2), ZN => l042_n_5);
  l042_g62 : CKAN2D1BWP7T port map(A1 => enable2, A2 => l042_n_3, Z => l042_n_4);
  l042_count_reg_0 : DFCNQD1BWP7T port map(CDN => l042_n_0, CP => clk, D => l042_n_2, Q => draw_count2(0));
  l042_g64 : CKXOR2D1BWP7T port map(A1 => draw_count2(0), A2 => draw_count2(1), Z => l042_n_3);
  l042_g65 : INR2XD0BWP7T port map(A1 => enable2, B1 => draw_count2(0), ZN => l042_n_2);
  l042_g66 : ND2D1BWP7T port map(A1 => draw_count2(1), A2 => draw_count2(0), ZN => l042_n_1);
  l042_g67 : INVD0BWP7T port map(I => reset, ZN => l042_n_0);
  l043_count_reg_2 : DFCNQD1BWP7T port map(CDN => l043_n_0, CP => clk, D => l043_n_6, Q => draw_count3(2));
  l043_g59 : CKAN2D1BWP7T port map(A1 => enable3, A2 => l043_n_5, Z => l043_n_6);
  l043_count_reg_1 : DFCNQD1BWP7T port map(CDN => l043_n_0, CP => clk, D => l043_n_4, Q => draw_count3(1));
  l043_g61 : MOAI22D0BWP7T port map(A1 => l043_n_1, A2 => draw_count3(2), B1 => l043_n_1, B2 => draw_count3(2), ZN => l043_n_5);
  l043_g62 : CKAN2D1BWP7T port map(A1 => enable3, A2 => l043_n_3, Z => l043_n_4);
  l043_count_reg_0 : DFCNQD1BWP7T port map(CDN => l043_n_0, CP => clk, D => l043_n_2, Q => draw_count3(0));
  l043_g64 : CKXOR2D1BWP7T port map(A1 => draw_count3(0), A2 => draw_count3(1), Z => l043_n_3);
  l043_g65 : INR2XD0BWP7T port map(A1 => enable3, B1 => draw_count3(0), ZN => l043_n_2);
  l043_g66 : ND2D1BWP7T port map(A1 => draw_count3(1), A2 => draw_count3(0), ZN => l043_n_1);
  l043_g67 : INVD0BWP7T port map(I => reset, ZN => l043_n_0);
  l044_count_reg_4 : DFCNQD1BWP7T port map(CDN => l044_n_0, CP => clk, D => l044_n_12, Q => draw_count4(4));
  l044_g82 : CKAN2D1BWP7T port map(A1 => enable4, A2 => l044_n_11, Z => l044_n_12);
  l044_count_reg_3 : DFCNQD1BWP7T port map(CDN => l044_n_0, CP => clk, D => l044_n_10, Q => draw_count4(3));
  l044_g84 : MOAI22D0BWP7T port map(A1 => l044_n_8, A2 => draw_count4(4), B1 => l044_n_8, B2 => draw_count4(4), ZN => l044_n_11);
  l044_g85 : CKAN2D1BWP7T port map(A1 => enable4, A2 => l044_n_9, Z => l044_n_10);
  l044_count_reg_2 : DFCNQD1BWP7T port map(CDN => l044_n_0, CP => clk, D => l044_n_7, Q => draw_count4(2));
  l044_g87 : MOAI22D0BWP7T port map(A1 => l044_n_4, A2 => draw_count4(3), B1 => l044_n_4, B2 => draw_count4(3), ZN => l044_n_9);
  l044_g88 : IND2D1BWP7T port map(A1 => l044_n_4, B1 => draw_count4(3), ZN => l044_n_8);
  l044_g89 : CKAN2D1BWP7T port map(A1 => enable4, A2 => l044_n_6, Z => l044_n_7);
  l044_count_reg_1 : DFCNQD1BWP7T port map(CDN => l044_n_0, CP => clk, D => l044_n_5, Q => draw_count4(1));
  l044_g91 : MOAI22D0BWP7T port map(A1 => l044_n_1, A2 => draw_count4(2), B1 => l044_n_1, B2 => draw_count4(2), ZN => l044_n_6);
  l044_g92 : CKAN2D1BWP7T port map(A1 => enable4, A2 => l044_n_3, Z => l044_n_5);
  l044_g93 : IND2D1BWP7T port map(A1 => l044_n_1, B1 => draw_count4(2), ZN => l044_n_4);
  l044_count_reg_0 : DFCNQD1BWP7T port map(CDN => l044_n_0, CP => clk, D => l044_n_2, Q => draw_count4(0));
  l044_g95 : CKXOR2D1BWP7T port map(A1 => draw_count4(0), A2 => draw_count4(1), Z => l044_n_3);
  l044_g96 : INR2XD0BWP7T port map(A1 => enable4, B1 => draw_count4(0), ZN => l044_n_2);
  l044_g97 : ND2D1BWP7T port map(A1 => draw_count4(1), A2 => draw_count4(0), ZN => l044_n_1);
  l044_g107 : INVD0BWP7T port map(I => reset, ZN => l044_n_0);
  l045_count_reg_4 : DFCNQD1BWP7T port map(CDN => l045_n_0, CP => clk, D => l045_n_12, Q => draw_count5(4));
  l045_g82 : CKAN2D1BWP7T port map(A1 => enable5, A2 => l045_n_11, Z => l045_n_12);
  l045_count_reg_3 : DFCNQD1BWP7T port map(CDN => l045_n_0, CP => clk, D => l045_n_10, Q => draw_count5(3));
  l045_g84 : MOAI22D0BWP7T port map(A1 => l045_n_8, A2 => draw_count5(4), B1 => l045_n_8, B2 => draw_count5(4), ZN => l045_n_11);
  l045_g85 : CKAN2D1BWP7T port map(A1 => enable5, A2 => l045_n_9, Z => l045_n_10);
  l045_count_reg_2 : DFCNQD1BWP7T port map(CDN => l045_n_0, CP => clk, D => l045_n_7, Q => draw_count5(2));
  l045_g87 : MOAI22D0BWP7T port map(A1 => l045_n_4, A2 => draw_count5(3), B1 => l045_n_4, B2 => draw_count5(3), ZN => l045_n_9);
  l045_g88 : IND2D1BWP7T port map(A1 => l045_n_4, B1 => draw_count5(3), ZN => l045_n_8);
  l045_g89 : CKAN2D1BWP7T port map(A1 => enable5, A2 => l045_n_6, Z => l045_n_7);
  l045_count_reg_1 : DFCNQD1BWP7T port map(CDN => l045_n_0, CP => clk, D => l045_n_5, Q => draw_count5(1));
  l045_g91 : MOAI22D0BWP7T port map(A1 => l045_n_1, A2 => draw_count5(2), B1 => l045_n_1, B2 => draw_count5(2), ZN => l045_n_6);
  l045_g92 : CKAN2D1BWP7T port map(A1 => enable5, A2 => l045_n_3, Z => l045_n_5);
  l045_g93 : IND2D1BWP7T port map(A1 => l045_n_1, B1 => draw_count5(2), ZN => l045_n_4);
  l045_count_reg_0 : DFCNQD1BWP7T port map(CDN => l045_n_0, CP => clk, D => l045_n_2, Q => draw_count5(0));
  l045_g95 : CKXOR2D1BWP7T port map(A1 => draw_count5(0), A2 => draw_count5(1), Z => l045_n_3);
  l045_g96 : INR2XD0BWP7T port map(A1 => enable5, B1 => draw_count5(0), ZN => l045_n_2);
  l045_g97 : ND2D1BWP7T port map(A1 => draw_count5(1), A2 => draw_count5(0), ZN => l045_n_1);
  l045_g107 : INVD0BWP7T port map(I => reset, ZN => l045_n_0);
  l046_count_reg_4 : DFCNQD1BWP7T port map(CDN => l046_n_0, CP => clk, D => l046_n_12, Q => draw_count6(4));
  l046_g82 : CKAN2D1BWP7T port map(A1 => enable6, A2 => l046_n_11, Z => l046_n_12);
  l046_count_reg_3 : DFCNQD1BWP7T port map(CDN => l046_n_0, CP => clk, D => l046_n_10, Q => draw_count6(3));
  l046_g84 : MOAI22D0BWP7T port map(A1 => l046_n_8, A2 => draw_count6(4), B1 => l046_n_8, B2 => draw_count6(4), ZN => l046_n_11);
  l046_g85 : CKAN2D1BWP7T port map(A1 => enable6, A2 => l046_n_9, Z => l046_n_10);
  l046_count_reg_2 : DFCNQD1BWP7T port map(CDN => l046_n_0, CP => clk, D => l046_n_7, Q => draw_count6(2));
  l046_g87 : MOAI22D0BWP7T port map(A1 => l046_n_4, A2 => draw_count6(3), B1 => l046_n_4, B2 => draw_count6(3), ZN => l046_n_9);
  l046_g88 : IND2D1BWP7T port map(A1 => l046_n_4, B1 => draw_count6(3), ZN => l046_n_8);
  l046_g89 : CKAN2D1BWP7T port map(A1 => enable6, A2 => l046_n_6, Z => l046_n_7);
  l046_count_reg_1 : DFCNQD1BWP7T port map(CDN => l046_n_0, CP => clk, D => l046_n_5, Q => draw_count6(1));
  l046_g91 : MOAI22D0BWP7T port map(A1 => l046_n_1, A2 => draw_count6(2), B1 => l046_n_1, B2 => draw_count6(2), ZN => l046_n_6);
  l046_g92 : CKAN2D1BWP7T port map(A1 => enable6, A2 => l046_n_3, Z => l046_n_5);
  l046_g93 : IND2D1BWP7T port map(A1 => l046_n_1, B1 => draw_count6(2), ZN => l046_n_4);
  l046_count_reg_0 : DFCNQD1BWP7T port map(CDN => l046_n_0, CP => clk, D => l046_n_2, Q => draw_count6(0));
  l046_g95 : CKXOR2D1BWP7T port map(A1 => draw_count6(0), A2 => draw_count6(1), Z => l046_n_3);
  l046_g96 : INR2XD0BWP7T port map(A1 => enable6, B1 => draw_count6(0), ZN => l046_n_2);
  l046_g97 : ND2D1BWP7T port map(A1 => draw_count6(1), A2 => draw_count6(0), ZN => l046_n_1);
  l046_g107 : INVD0BWP7T port map(I => reset, ZN => l046_n_0);
  l047_count_reg_4 : DFCNQD1BWP7T port map(CDN => l047_n_0, CP => clk, D => l047_n_12, Q => draw_count7(4));
  l047_g82 : CKAN2D1BWP7T port map(A1 => enable7, A2 => l047_n_11, Z => l047_n_12);
  l047_count_reg_3 : DFCNQD1BWP7T port map(CDN => l047_n_0, CP => clk, D => l047_n_10, Q => draw_count7(3));
  l047_g84 : MOAI22D0BWP7T port map(A1 => l047_n_8, A2 => draw_count7(4), B1 => l047_n_8, B2 => draw_count7(4), ZN => l047_n_11);
  l047_g85 : CKAN2D1BWP7T port map(A1 => enable7, A2 => l047_n_9, Z => l047_n_10);
  l047_count_reg_2 : DFCNQD1BWP7T port map(CDN => l047_n_0, CP => clk, D => l047_n_7, Q => draw_count7(2));
  l047_g87 : MOAI22D0BWP7T port map(A1 => l047_n_4, A2 => draw_count7(3), B1 => l047_n_4, B2 => draw_count7(3), ZN => l047_n_9);
  l047_g88 : IND2D1BWP7T port map(A1 => l047_n_4, B1 => draw_count7(3), ZN => l047_n_8);
  l047_g89 : CKAN2D1BWP7T port map(A1 => enable7, A2 => l047_n_6, Z => l047_n_7);
  l047_count_reg_1 : DFCNQD1BWP7T port map(CDN => l047_n_0, CP => clk, D => l047_n_5, Q => draw_count7(1));
  l047_g91 : MOAI22D0BWP7T port map(A1 => l047_n_1, A2 => draw_count7(2), B1 => l047_n_1, B2 => draw_count7(2), ZN => l047_n_6);
  l047_g92 : CKAN2D1BWP7T port map(A1 => enable7, A2 => l047_n_3, Z => l047_n_5);
  l047_g93 : IND2D1BWP7T port map(A1 => l047_n_1, B1 => draw_count7(2), ZN => l047_n_4);
  l047_count_reg_0 : DFCNQD1BWP7T port map(CDN => l047_n_0, CP => clk, D => l047_n_2, Q => draw_count7(0));
  l047_g95 : CKXOR2D1BWP7T port map(A1 => draw_count7(0), A2 => draw_count7(1), Z => l047_n_3);
  l047_g96 : INR2XD0BWP7T port map(A1 => enable7, B1 => draw_count7(0), ZN => l047_n_2);
  l047_g97 : ND2D1BWP7T port map(A1 => draw_count7(1), A2 => draw_count7(0), ZN => l047_n_1);
  l047_g107 : INVD0BWP7T port map(I => reset, ZN => l047_n_0);
  l048_count_reg_4 : DFCNQD1BWP7T port map(CDN => l048_n_0, CP => clk, D => l048_n_12, Q => draw_count8(4));
  l048_g82 : CKAN2D1BWP7T port map(A1 => enable8, A2 => l048_n_11, Z => l048_n_12);
  l048_count_reg_3 : DFCNQD1BWP7T port map(CDN => l048_n_0, CP => clk, D => l048_n_10, Q => draw_count8(3));
  l048_g84 : MOAI22D0BWP7T port map(A1 => l048_n_8, A2 => draw_count8(4), B1 => l048_n_8, B2 => draw_count8(4), ZN => l048_n_11);
  l048_g85 : CKAN2D1BWP7T port map(A1 => enable8, A2 => l048_n_9, Z => l048_n_10);
  l048_count_reg_2 : DFCNQD1BWP7T port map(CDN => l048_n_0, CP => clk, D => l048_n_7, Q => draw_count8(2));
  l048_g87 : MOAI22D0BWP7T port map(A1 => l048_n_4, A2 => draw_count8(3), B1 => l048_n_4, B2 => draw_count8(3), ZN => l048_n_9);
  l048_g88 : IND2D1BWP7T port map(A1 => l048_n_4, B1 => draw_count8(3), ZN => l048_n_8);
  l048_g89 : CKAN2D1BWP7T port map(A1 => enable8, A2 => l048_n_6, Z => l048_n_7);
  l048_count_reg_1 : DFCNQD1BWP7T port map(CDN => l048_n_0, CP => clk, D => l048_n_5, Q => draw_count8(1));
  l048_g91 : MOAI22D0BWP7T port map(A1 => l048_n_1, A2 => draw_count8(2), B1 => l048_n_1, B2 => draw_count8(2), ZN => l048_n_6);
  l048_g92 : CKAN2D1BWP7T port map(A1 => enable8, A2 => l048_n_3, Z => l048_n_5);
  l048_g93 : IND2D1BWP7T port map(A1 => l048_n_1, B1 => draw_count8(2), ZN => l048_n_4);
  l048_count_reg_0 : DFCNQD1BWP7T port map(CDN => l048_n_0, CP => clk, D => l048_n_2, Q => draw_count8(0));
  l048_g95 : CKXOR2D1BWP7T port map(A1 => draw_count8(0), A2 => draw_count8(1), Z => l048_n_3);
  l048_g96 : INR2XD0BWP7T port map(A1 => enable8, B1 => draw_count8(0), ZN => l048_n_2);
  l048_g97 : ND2D1BWP7T port map(A1 => draw_count8(1), A2 => draw_count8(0), ZN => l048_n_1);
  l048_g107 : INVD0BWP7T port map(I => reset, ZN => l048_n_0);
  l0410_count_reg_4 : DFCNQD1BWP7T port map(CDN => l0410_n_0, CP => clk, D => l0410_n_12, Q => draw_count10(4));
  l0410_g82 : CKAN2D1BWP7T port map(A1 => enable10, A2 => l0410_n_11, Z => l0410_n_12);
  l0410_count_reg_3 : DFCNQD1BWP7T port map(CDN => l0410_n_0, CP => clk, D => l0410_n_10, Q => draw_count10(3));
  l0410_g84 : MOAI22D0BWP7T port map(A1 => l0410_n_8, A2 => draw_count10(4), B1 => l0410_n_8, B2 => draw_count10(4), ZN => l0410_n_11);
  l0410_g85 : CKAN2D1BWP7T port map(A1 => enable10, A2 => l0410_n_9, Z => l0410_n_10);
  l0410_count_reg_2 : DFCNQD1BWP7T port map(CDN => l0410_n_0, CP => clk, D => l0410_n_7, Q => draw_count10(2));
  l0410_g87 : MOAI22D0BWP7T port map(A1 => l0410_n_4, A2 => draw_count10(3), B1 => l0410_n_4, B2 => draw_count10(3), ZN => l0410_n_9);
  l0410_g88 : IND2D1BWP7T port map(A1 => l0410_n_4, B1 => draw_count10(3), ZN => l0410_n_8);
  l0410_g89 : CKAN2D1BWP7T port map(A1 => enable10, A2 => l0410_n_6, Z => l0410_n_7);
  l0410_count_reg_1 : DFCNQD1BWP7T port map(CDN => l0410_n_0, CP => clk, D => l0410_n_5, Q => draw_count10(1));
  l0410_g91 : MOAI22D0BWP7T port map(A1 => l0410_n_1, A2 => draw_count10(2), B1 => l0410_n_1, B2 => draw_count10(2), ZN => l0410_n_6);
  l0410_g92 : CKAN2D1BWP7T port map(A1 => enable10, A2 => l0410_n_3, Z => l0410_n_5);
  l0410_g93 : IND2D1BWP7T port map(A1 => l0410_n_1, B1 => draw_count10(2), ZN => l0410_n_4);
  l0410_count_reg_0 : DFCNQD1BWP7T port map(CDN => l0410_n_0, CP => clk, D => l0410_n_2, Q => draw_count10(0));
  l0410_g95 : CKXOR2D1BWP7T port map(A1 => draw_count10(0), A2 => draw_count10(1), Z => l0410_n_3);
  l0410_g96 : INR2XD0BWP7T port map(A1 => enable10, B1 => draw_count10(0), ZN => l0410_n_2);
  l0410_g97 : ND2D1BWP7T port map(A1 => draw_count10(1), A2 => draw_count10(0), ZN => l0410_n_1);
  l0410_g107 : INVD0BWP7T port map(I => reset, ZN => l0410_n_0);
  l049_count_reg_4 : DFCNQD1BWP7T port map(CDN => l049_n_0, CP => clk, D => l049_n_12, Q => draw_count9(4));
  l049_g82 : CKAN2D1BWP7T port map(A1 => enable9, A2 => l049_n_11, Z => l049_n_12);
  l049_count_reg_3 : DFCNQD1BWP7T port map(CDN => l049_n_0, CP => clk, D => l049_n_10, Q => draw_count9(3));
  l049_g84 : MOAI22D0BWP7T port map(A1 => l049_n_8, A2 => draw_count9(4), B1 => l049_n_8, B2 => draw_count9(4), ZN => l049_n_11);
  l049_g85 : CKAN2D1BWP7T port map(A1 => enable9, A2 => l049_n_9, Z => l049_n_10);
  l049_count_reg_2 : DFCNQD1BWP7T port map(CDN => l049_n_0, CP => clk, D => l049_n_7, Q => draw_count9(2));
  l049_g87 : MOAI22D0BWP7T port map(A1 => l049_n_4, A2 => draw_count9(3), B1 => l049_n_4, B2 => draw_count9(3), ZN => l049_n_9);
  l049_g88 : IND2D1BWP7T port map(A1 => l049_n_4, B1 => draw_count9(3), ZN => l049_n_8);
  l049_g89 : CKAN2D1BWP7T port map(A1 => enable9, A2 => l049_n_6, Z => l049_n_7);
  l049_count_reg_1 : DFCNQD1BWP7T port map(CDN => l049_n_0, CP => clk, D => l049_n_5, Q => draw_count9(1));
  l049_g91 : MOAI22D0BWP7T port map(A1 => l049_n_1, A2 => draw_count9(2), B1 => l049_n_1, B2 => draw_count9(2), ZN => l049_n_6);
  l049_g92 : CKAN2D1BWP7T port map(A1 => enable9, A2 => l049_n_3, Z => l049_n_5);
  l049_g93 : IND2D1BWP7T port map(A1 => l049_n_1, B1 => draw_count9(2), ZN => l049_n_4);
  l049_count_reg_0 : DFCNQD1BWP7T port map(CDN => l049_n_0, CP => clk, D => l049_n_2, Q => draw_count9(0));
  l049_g95 : CKXOR2D1BWP7T port map(A1 => draw_count9(0), A2 => draw_count9(1), Z => l049_n_3);
  l049_g96 : INR2XD0BWP7T port map(A1 => enable9, B1 => draw_count9(0), ZN => l049_n_2);
  l049_g97 : ND2D1BWP7T port map(A1 => draw_count9(1), A2 => draw_count9(0), ZN => l049_n_1);
  l049_g107 : INVD0BWP7T port map(I => reset, ZN => l049_n_0);
  l051_g2484 : OA21D0BWP7T port map(A1 => l051_n_82, A2 => l051_n_39, B => enable1, Z => r1);
  l051_g2485 : AO31D1BWP7T port map(A1 => l051_n_79, A2 => l051_n_77, A3 => draw_count1(0), B => b1, Z => g1);
  l051_g2486 : AO31D1BWP7T port map(A1 => l051_n_79, A2 => l051_n_77, A3 => l051_n_15, B => l051_n_83, Z => b1);
  l051_g2487 : OA21D0BWP7T port map(A1 => l051_n_80, A2 => l051_n_78, B => l051_n_39, Z => l051_n_83);
  l051_g2488 : OAI22D0BWP7T port map(A1 => l051_n_80, A2 => l051_n_73, B1 => l051_n_2, B2 => draw_count1(2), ZN => l051_n_82);
  l051_g2489 : OR2D1BWP7T port map(A1 => l051_n_77, A2 => l051_n_78, Z => enable1);
  l051_g2490 : INVD0BWP7T port map(I => l051_n_80, ZN => l051_n_79);
  l051_g2491 : NR2D1BWP7T port map(A1 => l051_n_76, A2 => l051_n_74, ZN => l051_n_80);
  l051_g2492 : INR2D1BWP7T port map(A1 => l051_n_73, B1 => l051_n_76, ZN => l051_n_78);
  l051_g2493 : AOI21D0BWP7T port map(A1 => l051_n_74, A2 => l051_n_0, B => l051_n_76, ZN => l051_n_77);
  l051_g2494 : OAI221D0BWP7T port map(A1 => l051_n_31, A2 => l051_n_9, B1 => l051_n_10, B2 => l051_n_33, C => l051_n_75, ZN => l051_n_76);
  l051_g2495 : NR4D0BWP7T port map(A1 => l051_n_71, A2 => l051_n_67, A3 => l051_n_60, A4 => l051_n_53, ZN => l051_n_75);
  l051_g2497 : ND4D0BWP7T port map(A1 => l051_n_72, A2 => l051_n_57, A3 => l051_n_35, A4 => l051_n_29, ZN => l051_n_74);
  l051_g2498 : NR4D0BWP7T port map(A1 => l051_n_70, A2 => l051_n_35, A3 => l051_n_36, A4 => l051_n_26, ZN => l051_n_73);
  l051_g2499 : AOI211XD0BWP7T port map(A1 => l051_n_30, A2 => l051_n_16, B => l051_n_69, C => l051_n_63, ZN => l051_n_72);
  l051_g2500 : OAI211D1BWP7T port map(A1 => l051_n_14, A2 => l051_n_25, B => l051_n_68, C => l051_n_51, ZN => l051_n_71);
  l051_g2501 : ND4D0BWP7T port map(A1 => l051_n_65, A2 => l051_n_61, A3 => l051_n_37, A4 => l051_n_29, ZN => l051_n_70);
  l051_g2502 : OAI211D1BWP7T port map(A1 => l051_n_16, A2 => l051_n_30, B => l051_n_66, C => l051_n_56, ZN => l051_n_69);
  l051_g2503 : MAOI222D1BWP7T port map(A => l051_n_64, B => l051_n_34, C => l051_n_5, ZN => l051_n_68);
  l051_g2504 : AOI22D0BWP7T port map(A1 => l051_n_62, A2 => l051_n_52, B1 => l051_n_34, B2 => l051_n_18, ZN => l051_n_67);
  l051_g2505 : AN3D1BWP7T port map(A1 => l051_n_55, A2 => l051_n_50, A3 => l051_n_61, Z => l051_n_66);
  l051_g2506 : NR3D0BWP7T port map(A1 => l051_n_63, A2 => l051_n_54, A3 => l051_n_30, ZN => l051_n_65);
  l051_g2507 : MAOI222D1BWP7T port map(A => l051_n_48, B => l051_n_28, C => x(2), ZN => l051_n_64);
  l051_g2508 : OAI211D1BWP7T port map(A1 => l051_n_17, A2 => l051_n_32, B => l051_n_47, C => l051_n_59, ZN => l051_n_63);
  l051_g2509 : AO211D0BWP7T port map(A1 => l051_n_28, A2 => l051_n_19, B => l051_n_46, C => l051_n_42, Z => l051_n_62);
  l051_g2510 : MOAI22D0BWP7T port map(A1 => x(8), A2 => l051_n_1, B1 => l051_n_31, B2 => l051_n_9, ZN => l051_n_60);
  l051_g2511 : MAOI22D0BWP7T port map(A1 => l051_n_20, A2 => y(9), B1 => l051_n_20, B2 => y(9), ZN => l051_n_59);
  l051_g2512 : MAOI22D0BWP7T port map(A1 => l051_n_26, A2 => l051_n_13, B1 => l051_n_26, B2 => l051_n_13, ZN => l051_n_58);
  l051_g2513 : MAOI22D0BWP7T port map(A1 => l051_n_26, A2 => y(1), B1 => l051_n_26, B2 => y(1), ZN => l051_n_57);
  l051_g2514 : MAOI22D0BWP7T port map(A1 => l051_n_37, A2 => l051_n_11, B1 => l051_n_37, B2 => l051_n_11, ZN => l051_n_56);
  l051_g2515 : MOAI22D0BWP7T port map(A1 => l051_n_38, A2 => l051_n_12, B1 => l051_n_38, B2 => l051_n_12, ZN => l051_n_61);
  l051_g2516 : MAOI22D0BWP7T port map(A1 => l051_n_45, A2 => l051_n_44, B1 => l051_n_36, B2 => l051_n_22, ZN => l051_n_55);
  l051_g2517 : MOAI22D0BWP7T port map(A1 => l051_n_45, A2 => y(5), B1 => l051_n_45, B2 => y(5), ZN => l051_n_54);
  l051_g2518 : MOAI22D0BWP7T port map(A1 => l051_n_40, A2 => l051_n_24, B1 => l051_n_14, B2 => l051_n_25, ZN => l051_n_53);
  l051_g2519 : OA22D0BWP7T port map(A1 => l051_n_34, A2 => l051_n_18, B1 => l051_n_19, B2 => l051_n_28, Z => l051_n_52);
  l051_g2520 : AOI22D0BWP7T port map(A1 => l051_n_40, A2 => l051_n_24, B1 => l051_n_33, B2 => l051_n_10, ZN => l051_n_51);
  l051_g2521 : AOI22D0BWP7T port map(A1 => l051_n_36, A2 => l051_n_22, B1 => l051_n_27, B2 => l051_n_7, ZN => l051_n_50);
  l051_g2522 : MAOI22D0BWP7T port map(A1 => l051_n_35, A2 => y(0), B1 => l051_n_35, B2 => y(0), ZN => l051_n_49);
  l051_g2523 : OR2D1BWP7T port map(A1 => l051_n_43, A2 => l051_n_6, Z => l051_n_48);
  l051_g2524 : ND2D1BWP7T port map(A1 => l051_n_32, A2 => l051_n_17, ZN => l051_n_47);
  l051_g2525 : OA21D0BWP7T port map(A1 => l051_n_41, A2 => l051_n_6, B => l051_n_23, Z => l051_n_46);
  l051_g2526 : INVD0BWP7T port map(I => l051_n_27, ZN => l051_n_45);
  l051_g2527 : INVD0BWP7T port map(I => l051_n_7, ZN => l051_n_44);
  l051_g2528 : AOI21D0BWP7T port map(A1 => l051_n_21, A2 => l051_n_23, B => l051_n_41, ZN => l051_n_43);
  l051_g2529 : OA21D0BWP7T port map(A1 => l051_n_8, A2 => l051_n_6, B => l051_n_21, Z => l051_n_42);
  l051_g2530 : AO21D0BWP7T port map(A1 => l051_n_4, A2 => x_bullet1(1), B => l051_n_8, Z => l051_n_41);
  l051_g2531 : MAOI22D0BWP7T port map(A1 => x(6), A2 => x_bullet1(6), B1 => x(6), B2 => x_bullet1(6), ZN => l051_n_40);
  l051_g2532 : OA21D0BWP7T port map(A1 => l051_n_2, A2 => draw_count1(1), B => l051_n_15, Z => l051_n_39);
  l051_g2533 : MOAI22D0BWP7T port map(A1 => y(7), A2 => y_bullet1(7), B1 => y(7), B2 => y_bullet1(7), ZN => l051_n_38);
  l051_g2534 : OAI21D0BWP7T port map(A1 => y(5), A2 => l051_n_3, B => l051_n_7, ZN => l051_n_37);
  l051_g2535 : MAOI22D0BWP7T port map(A1 => y(4), A2 => y_bullet1(4), B1 => y(4), B2 => y_bullet1(4), ZN => l051_n_36);
  l051_g2536 : MAOI22D0BWP7T port map(A1 => y(1), A2 => y_bullet1(1), B1 => y(1), B2 => y_bullet1(1), ZN => l051_n_35);
  l051_g2537 : MOAI22D0BWP7T port map(A1 => x(4), A2 => x_bullet1(4), B1 => x(4), B2 => x_bullet1(4), ZN => l051_n_34);
  l051_g2539 : MOAI22D0BWP7T port map(A1 => x(5), A2 => x_bullet1(5), B1 => x(5), B2 => x_bullet1(5), ZN => l051_n_33);
  l051_g2540 : MOAI22D0BWP7T port map(A1 => y(8), A2 => y_bullet1(8), B1 => y(8), B2 => y_bullet1(8), ZN => l051_n_32);
  l051_g2541 : MOAI22D0BWP7T port map(A1 => x(7), A2 => x_bullet1(7), B1 => x(7), B2 => x_bullet1(7), ZN => l051_n_31);
  l051_g2542 : MAOI22D0BWP7T port map(A1 => y(3), A2 => y_bullet1(3), B1 => y(3), B2 => y_bullet1(3), ZN => l051_n_30);
  l051_g2543 : MOAI22D0BWP7T port map(A1 => y(0), A2 => y_bullet1(0), B1 => y(0), B2 => y_bullet1(0), ZN => l051_n_29);
  l051_g2544 : MAOI22D0BWP7T port map(A1 => x(3), A2 => x_bullet1(3), B1 => x(3), B2 => x_bullet1(3), ZN => l051_n_28);
  l051_g2545 : MOAI22D0BWP7T port map(A1 => y(6), A2 => y_bullet1(6), B1 => y(6), B2 => y_bullet1(6), ZN => l051_n_27);
  l051_g2546 : MAOI22D0BWP7T port map(A1 => y(2), A2 => y_bullet1(2), B1 => y(2), B2 => y_bullet1(2), ZN => l051_n_26);
  l051_g2547 : IND2D1BWP7T port map(A1 => x(7), B1 => x_bullet1(7), ZN => l051_n_25);
  l051_g2548 : INR2D0BWP7T port map(A1 => x_bullet1(5), B1 => x(5), ZN => l051_n_24);
  l051_g2549 : IND2D0BWP7T port map(A1 => x_bullet1(0), B1 => x(0), ZN => l051_n_23);
  l051_g2550 : IND2D1BWP7T port map(A1 => y(3), B1 => y_bullet1(3), ZN => l051_n_22);
  l051_g2551 : IND2D0BWP7T port map(A1 => x_bullet1(1), B1 => x(1), ZN => l051_n_21);
  l051_g2552 : IND2D1BWP7T port map(A1 => y(8), B1 => y_bullet1(8), ZN => l051_n_20);
  l051_g2553 : INR2D0BWP7T port map(A1 => x_bullet1(2), B1 => x(2), ZN => l051_n_19);
  l051_g2554 : IND2D0BWP7T port map(A1 => x_bullet1(3), B1 => x(3), ZN => l051_n_18);
  l051_g2555 : INR2XD0BWP7T port map(A1 => y_bullet1(7), B1 => y(7), ZN => l051_n_17);
  l051_g2556 : IND2D1BWP7T port map(A1 => y(2), B1 => y_bullet1(2), ZN => l051_n_16);
  l051_g2557 : OR2D1BWP7T port map(A1 => draw_count1(1), A2 => draw_count1(2), Z => l051_n_15);
  l051_g2558 : AN2D1BWP7T port map(A1 => x(8), A2 => l051_n_1, Z => l051_n_14);
  l051_g2559 : INR2D0BWP7T port map(A1 => x_bullet1(3), B1 => x(3), ZN => l051_n_5);
  l051_g2560 : IND2D1BWP7T port map(A1 => y(1), B1 => y_bullet1(1), ZN => l051_n_13);
  l051_g2561 : IND2D1BWP7T port map(A1 => y(6), B1 => y_bullet1(6), ZN => l051_n_12);
  l051_g2562 : INR2XD0BWP7T port map(A1 => y_bullet1(4), B1 => y(4), ZN => l051_n_11);
  l051_g2563 : INR2D0BWP7T port map(A1 => x_bullet1(4), B1 => x(4), ZN => l051_n_10);
  l051_g2564 : IND2D0BWP7T port map(A1 => x_bullet1(6), B1 => x(6), ZN => l051_n_9);
  l051_g2565 : AN2D0BWP7T port map(A1 => x(2), A2 => x_bullet1(2), Z => l051_n_8);
  l051_g2566 : ND2D1BWP7T port map(A1 => y(5), A2 => l051_n_3, ZN => l051_n_7);
  l051_g2567 : NR2D0BWP7T port map(A1 => x(2), A2 => x_bullet1(2), ZN => l051_n_6);
  l051_g2568 : INVD0BWP7T port map(I => x(1), ZN => l051_n_4);
  l051_g2569 : INVD1BWP7T port map(I => y_bullet1(5), ZN => l051_n_3);
  l051_g2570 : INVD0BWP7T port map(I => draw_count1(0), ZN => l051_n_2);
  l051_g2571 : INVD0BWP7T port map(I => x_bullet1(8), ZN => l051_n_1);
  l051_g2 : IND4D0BWP7T port map(A1 => l051_n_29, B1 => l051_n_72, B2 => l051_n_49, B3 => l051_n_58, ZN => l051_n_0);
  l052_g2484 : OA21D0BWP7T port map(A1 => l052_n_82, A2 => l052_n_39, B => enable2, Z => r2);
  l052_g2485 : AO31D1BWP7T port map(A1 => l052_n_79, A2 => l052_n_77, A3 => draw_count2(0), B => b2, Z => g2);
  l052_g2486 : AO31D1BWP7T port map(A1 => l052_n_79, A2 => l052_n_77, A3 => l052_n_15, B => l052_n_83, Z => b2);
  l052_g2487 : OA21D0BWP7T port map(A1 => l052_n_80, A2 => l052_n_78, B => l052_n_39, Z => l052_n_83);
  l052_g2488 : OAI22D0BWP7T port map(A1 => l052_n_80, A2 => l052_n_73, B1 => l052_n_2, B2 => draw_count2(2), ZN => l052_n_82);
  l052_g2489 : OR2D1BWP7T port map(A1 => l052_n_77, A2 => l052_n_78, Z => enable2);
  l052_g2490 : INVD0BWP7T port map(I => l052_n_80, ZN => l052_n_79);
  l052_g2491 : NR2D1BWP7T port map(A1 => l052_n_76, A2 => l052_n_74, ZN => l052_n_80);
  l052_g2492 : INR2D1BWP7T port map(A1 => l052_n_73, B1 => l052_n_76, ZN => l052_n_78);
  l052_g2493 : AOI21D0BWP7T port map(A1 => l052_n_74, A2 => l052_n_0, B => l052_n_76, ZN => l052_n_77);
  l052_g2494 : OAI221D0BWP7T port map(A1 => l052_n_31, A2 => l052_n_9, B1 => l052_n_10, B2 => l052_n_33, C => l052_n_75, ZN => l052_n_76);
  l052_g2495 : NR4D0BWP7T port map(A1 => l052_n_71, A2 => l052_n_67, A3 => l052_n_60, A4 => l052_n_53, ZN => l052_n_75);
  l052_g2497 : ND4D0BWP7T port map(A1 => l052_n_72, A2 => l052_n_57, A3 => l052_n_35, A4 => l052_n_29, ZN => l052_n_74);
  l052_g2498 : NR4D0BWP7T port map(A1 => l052_n_70, A2 => l052_n_35, A3 => l052_n_36, A4 => l052_n_26, ZN => l052_n_73);
  l052_g2499 : AOI211XD0BWP7T port map(A1 => l052_n_30, A2 => l052_n_16, B => l052_n_69, C => l052_n_63, ZN => l052_n_72);
  l052_g2500 : OAI211D1BWP7T port map(A1 => l052_n_14, A2 => l052_n_25, B => l052_n_68, C => l052_n_51, ZN => l052_n_71);
  l052_g2501 : ND4D0BWP7T port map(A1 => l052_n_65, A2 => l052_n_61, A3 => l052_n_37, A4 => l052_n_29, ZN => l052_n_70);
  l052_g2502 : OAI211D1BWP7T port map(A1 => l052_n_16, A2 => l052_n_30, B => l052_n_66, C => l052_n_56, ZN => l052_n_69);
  l052_g2503 : MAOI222D1BWP7T port map(A => l052_n_64, B => l052_n_34, C => l052_n_5, ZN => l052_n_68);
  l052_g2504 : AOI22D0BWP7T port map(A1 => l052_n_62, A2 => l052_n_52, B1 => l052_n_34, B2 => l052_n_18, ZN => l052_n_67);
  l052_g2505 : AN3D1BWP7T port map(A1 => l052_n_55, A2 => l052_n_50, A3 => l052_n_61, Z => l052_n_66);
  l052_g2506 : NR3D0BWP7T port map(A1 => l052_n_63, A2 => l052_n_54, A3 => l052_n_30, ZN => l052_n_65);
  l052_g2507 : MAOI222D1BWP7T port map(A => l052_n_48, B => l052_n_28, C => x(2), ZN => l052_n_64);
  l052_g2508 : OAI211D1BWP7T port map(A1 => l052_n_17, A2 => l052_n_32, B => l052_n_47, C => l052_n_59, ZN => l052_n_63);
  l052_g2509 : AO211D0BWP7T port map(A1 => l052_n_28, A2 => l052_n_19, B => l052_n_46, C => l052_n_42, Z => l052_n_62);
  l052_g2510 : MOAI22D0BWP7T port map(A1 => x(8), A2 => l052_n_1, B1 => l052_n_31, B2 => l052_n_9, ZN => l052_n_60);
  l052_g2511 : MAOI22D0BWP7T port map(A1 => l052_n_20, A2 => y(9), B1 => l052_n_20, B2 => y(9), ZN => l052_n_59);
  l052_g2512 : MAOI22D0BWP7T port map(A1 => l052_n_26, A2 => l052_n_13, B1 => l052_n_26, B2 => l052_n_13, ZN => l052_n_58);
  l052_g2513 : MAOI22D0BWP7T port map(A1 => l052_n_26, A2 => y(1), B1 => l052_n_26, B2 => y(1), ZN => l052_n_57);
  l052_g2514 : MAOI22D0BWP7T port map(A1 => l052_n_37, A2 => l052_n_11, B1 => l052_n_37, B2 => l052_n_11, ZN => l052_n_56);
  l052_g2515 : MOAI22D0BWP7T port map(A1 => l052_n_38, A2 => l052_n_12, B1 => l052_n_38, B2 => l052_n_12, ZN => l052_n_61);
  l052_g2516 : MAOI22D0BWP7T port map(A1 => l052_n_45, A2 => l052_n_44, B1 => l052_n_36, B2 => l052_n_22, ZN => l052_n_55);
  l052_g2517 : MOAI22D0BWP7T port map(A1 => l052_n_45, A2 => y(5), B1 => l052_n_45, B2 => y(5), ZN => l052_n_54);
  l052_g2518 : MOAI22D0BWP7T port map(A1 => l052_n_40, A2 => l052_n_24, B1 => l052_n_14, B2 => l052_n_25, ZN => l052_n_53);
  l052_g2519 : OA22D0BWP7T port map(A1 => l052_n_34, A2 => l052_n_18, B1 => l052_n_19, B2 => l052_n_28, Z => l052_n_52);
  l052_g2520 : AOI22D0BWP7T port map(A1 => l052_n_40, A2 => l052_n_24, B1 => l052_n_33, B2 => l052_n_10, ZN => l052_n_51);
  l052_g2521 : AOI22D0BWP7T port map(A1 => l052_n_36, A2 => l052_n_22, B1 => l052_n_27, B2 => l052_n_7, ZN => l052_n_50);
  l052_g2522 : MAOI22D0BWP7T port map(A1 => l052_n_35, A2 => y(0), B1 => l052_n_35, B2 => y(0), ZN => l052_n_49);
  l052_g2523 : OR2D1BWP7T port map(A1 => l052_n_43, A2 => l052_n_6, Z => l052_n_48);
  l052_g2524 : ND2D1BWP7T port map(A1 => l052_n_32, A2 => l052_n_17, ZN => l052_n_47);
  l052_g2525 : OA21D0BWP7T port map(A1 => l052_n_41, A2 => l052_n_6, B => l052_n_23, Z => l052_n_46);
  l052_g2526 : INVD0BWP7T port map(I => l052_n_27, ZN => l052_n_45);
  l052_g2527 : INVD0BWP7T port map(I => l052_n_7, ZN => l052_n_44);
  l052_g2528 : AOI21D0BWP7T port map(A1 => l052_n_21, A2 => l052_n_23, B => l052_n_41, ZN => l052_n_43);
  l052_g2529 : OA21D0BWP7T port map(A1 => l052_n_8, A2 => l052_n_6, B => l052_n_21, Z => l052_n_42);
  l052_g2530 : AO21D0BWP7T port map(A1 => l052_n_4, A2 => x_bullet2(1), B => l052_n_8, Z => l052_n_41);
  l052_g2531 : MAOI22D0BWP7T port map(A1 => x(6), A2 => x_bullet2(6), B1 => x(6), B2 => x_bullet2(6), ZN => l052_n_40);
  l052_g2532 : OA21D0BWP7T port map(A1 => l052_n_2, A2 => draw_count2(1), B => l052_n_15, Z => l052_n_39);
  l052_g2533 : MOAI22D0BWP7T port map(A1 => y(7), A2 => y_bullet2(7), B1 => y(7), B2 => y_bullet2(7), ZN => l052_n_38);
  l052_g2534 : OAI21D0BWP7T port map(A1 => y(5), A2 => l052_n_3, B => l052_n_7, ZN => l052_n_37);
  l052_g2535 : MAOI22D0BWP7T port map(A1 => y(4), A2 => y_bullet2(4), B1 => y(4), B2 => y_bullet2(4), ZN => l052_n_36);
  l052_g2536 : MAOI22D0BWP7T port map(A1 => y(1), A2 => y_bullet2(1), B1 => y(1), B2 => y_bullet2(1), ZN => l052_n_35);
  l052_g2537 : MOAI22D0BWP7T port map(A1 => x(4), A2 => x_bullet2(4), B1 => x(4), B2 => x_bullet2(4), ZN => l052_n_34);
  l052_g2539 : MOAI22D0BWP7T port map(A1 => x(5), A2 => x_bullet2(5), B1 => x(5), B2 => x_bullet2(5), ZN => l052_n_33);
  l052_g2540 : MOAI22D0BWP7T port map(A1 => y(8), A2 => y_bullet2(8), B1 => y(8), B2 => y_bullet2(8), ZN => l052_n_32);
  l052_g2541 : MOAI22D0BWP7T port map(A1 => x(7), A2 => x_bullet2(7), B1 => x(7), B2 => x_bullet2(7), ZN => l052_n_31);
  l052_g2542 : MAOI22D0BWP7T port map(A1 => y(3), A2 => y_bullet2(3), B1 => y(3), B2 => y_bullet2(3), ZN => l052_n_30);
  l052_g2543 : MOAI22D0BWP7T port map(A1 => y(0), A2 => y_bullet2(0), B1 => y(0), B2 => y_bullet2(0), ZN => l052_n_29);
  l052_g2544 : MAOI22D0BWP7T port map(A1 => x(3), A2 => x_bullet2(3), B1 => x(3), B2 => x_bullet2(3), ZN => l052_n_28);
  l052_g2545 : MOAI22D0BWP7T port map(A1 => y(6), A2 => y_bullet2(6), B1 => y(6), B2 => y_bullet2(6), ZN => l052_n_27);
  l052_g2546 : MAOI22D0BWP7T port map(A1 => y(2), A2 => y_bullet2(2), B1 => y(2), B2 => y_bullet2(2), ZN => l052_n_26);
  l052_g2547 : IND2D1BWP7T port map(A1 => x(7), B1 => x_bullet2(7), ZN => l052_n_25);
  l052_g2548 : INR2D0BWP7T port map(A1 => x_bullet2(5), B1 => x(5), ZN => l052_n_24);
  l052_g2549 : IND2D0BWP7T port map(A1 => x_bullet2(0), B1 => x(0), ZN => l052_n_23);
  l052_g2550 : IND2D1BWP7T port map(A1 => y(3), B1 => y_bullet2(3), ZN => l052_n_22);
  l052_g2551 : IND2D0BWP7T port map(A1 => x_bullet2(1), B1 => x(1), ZN => l052_n_21);
  l052_g2552 : IND2D1BWP7T port map(A1 => y(8), B1 => y_bullet2(8), ZN => l052_n_20);
  l052_g2553 : INR2D0BWP7T port map(A1 => x_bullet2(2), B1 => x(2), ZN => l052_n_19);
  l052_g2554 : IND2D0BWP7T port map(A1 => x_bullet2(3), B1 => x(3), ZN => l052_n_18);
  l052_g2555 : INR2XD0BWP7T port map(A1 => y_bullet2(7), B1 => y(7), ZN => l052_n_17);
  l052_g2556 : IND2D1BWP7T port map(A1 => y(2), B1 => y_bullet2(2), ZN => l052_n_16);
  l052_g2557 : OR2D1BWP7T port map(A1 => draw_count2(1), A2 => draw_count2(2), Z => l052_n_15);
  l052_g2558 : AN2D1BWP7T port map(A1 => x(8), A2 => l052_n_1, Z => l052_n_14);
  l052_g2559 : INR2D0BWP7T port map(A1 => x_bullet2(3), B1 => x(3), ZN => l052_n_5);
  l052_g2560 : IND2D1BWP7T port map(A1 => y(1), B1 => y_bullet2(1), ZN => l052_n_13);
  l052_g2561 : IND2D1BWP7T port map(A1 => y(6), B1 => y_bullet2(6), ZN => l052_n_12);
  l052_g2562 : INR2XD0BWP7T port map(A1 => y_bullet2(4), B1 => y(4), ZN => l052_n_11);
  l052_g2563 : INR2D0BWP7T port map(A1 => x_bullet2(4), B1 => x(4), ZN => l052_n_10);
  l052_g2564 : IND2D0BWP7T port map(A1 => x_bullet2(6), B1 => x(6), ZN => l052_n_9);
  l052_g2565 : AN2D0BWP7T port map(A1 => x(2), A2 => x_bullet2(2), Z => l052_n_8);
  l052_g2566 : ND2D1BWP7T port map(A1 => y(5), A2 => l052_n_3, ZN => l052_n_7);
  l052_g2567 : NR2D0BWP7T port map(A1 => x(2), A2 => x_bullet2(2), ZN => l052_n_6);
  l052_g2568 : INVD0BWP7T port map(I => x(1), ZN => l052_n_4);
  l052_g2569 : INVD1BWP7T port map(I => y_bullet2(5), ZN => l052_n_3);
  l052_g2570 : INVD0BWP7T port map(I => draw_count2(0), ZN => l052_n_2);
  l052_g2571 : INVD0BWP7T port map(I => x_bullet2(8), ZN => l052_n_1);
  l052_g2 : IND4D0BWP7T port map(A1 => l052_n_29, B1 => l052_n_72, B2 => l052_n_49, B3 => l052_n_58, ZN => l052_n_0);
  l071_g12395 : OAI221D0BWP7T port map(A1 => l071_n_222, A2 => l071_n_184, B1 => l071_n_156, B2 => l071_n_225, C => l071_n_246, ZN => r5);
  l071_g12396 : NR4D0BWP7T port map(A1 => l071_n_245, A2 => l071_n_235, A3 => l071_n_229, A4 => l071_n_206, ZN => l071_n_246);
  l071_g12397 : IND4D0BWP7T port map(A1 => l071_n_233, B1 => l071_n_228, B2 => l071_n_234, B3 => l071_n_242, ZN => l071_n_245);
  l071_g12398 : AO211D0BWP7T port map(A1 => l071_n_218, A2 => l071_n_92, B => l071_n_243, C => l071_n_241, Z => g5);
  l071_g12399 : OAI211D1BWP7T port map(A1 => l071_n_126, A2 => l071_n_222, B => l071_n_239, C => l071_n_231, ZN => l071_n_243);
  l071_g12400 : MAOI22D0BWP7T port map(A1 => l071_n_215, A2 => l071_n_162, B1 => l071_n_236, B2 => l071_n_194, ZN => l071_n_242);
  l071_g12401 : AO221D0BWP7T port map(A1 => l071_n_215, A2 => l071_n_139, B1 => l071_n_212, B2 => l071_n_127, C => l071_n_237, Z => l071_n_241);
  l071_g12402 : OAI32D1BWP7T port map(A1 => l071_n_25, A2 => l071_n_61, A3 => l071_n_222, B1 => l071_n_96, B2 => l071_n_224, ZN => b5);
  l071_g12403 : AOI211XD0BWP7T port map(A1 => l071_n_199, A2 => l071_n_71, B => l071_n_232, C => l071_n_226, ZN => l071_n_239);
  l071_g12404 : ND3D0BWP7T port map(A1 => l071_n_220, A2 => l071_n_211, A3 => l071_n_198, ZN => enable5);
  l071_g12405 : OAI211D1BWP7T port map(A1 => l071_n_85, A2 => l071_n_204, B => l071_n_219, C => l071_n_227, ZN => l071_n_237);
  l071_g12406 : ND4D0BWP7T port map(A1 => l071_n_216, A2 => l071_n_187, A3 => l071_n_181, A4 => l071_n_165, ZN => l071_n_236);
  l071_g12407 : OAI211D1BWP7T port map(A1 => l071_n_172, A2 => l071_n_224, B => l071_n_221, C => l071_n_207, ZN => l071_n_235);
  l071_g12408 : AOI22D0BWP7T port map(A1 => l071_n_212, A2 => l071_n_157, B1 => l071_n_217, B2 => l071_n_161, ZN => l071_n_234);
  l071_g12409 : AOI31D0BWP7T port map(A1 => l071_n_132, A2 => l071_n_130, A3 => l071_n_61, B => l071_n_230, ZN => l071_n_233);
  l071_g12410 : AOI21D0BWP7T port map(A1 => l071_n_132, A2 => l071_n_72, B => l071_n_225, ZN => l071_n_232);
  l071_g12411 : OAI21D0BWP7T port map(A1 => l071_n_133, A2 => l071_n_92, B => l071_n_223, ZN => l071_n_231);
  l071_g12412 : AOI21D0BWP7T port map(A1 => l071_n_210, A2 => l071_n_150, B => l071_n_196, ZN => l071_n_230);
  l071_g12413 : IAO21D0BWP7T port map(A1 => l071_n_153, A2 => l071_n_71, B => l071_n_213, ZN => l071_n_229);
  l071_g12414 : OAI31D0BWP7T port map(A1 => l071_n_76, A2 => l071_n_112, A3 => l071_n_92, B => l071_n_214, ZN => l071_n_228);
  l071_g12415 : OAI21D0BWP7T port map(A1 => l071_n_133, A2 => l071_n_139, B => l071_n_214, ZN => l071_n_227);
  l071_g12416 : AOI21D0BWP7T port map(A1 => l071_n_103, A2 => l071_n_70, B => l071_n_213, ZN => l071_n_226);
  l071_g12417 : INVD0BWP7T port map(I => l071_n_223, ZN => l071_n_224);
  l071_g12418 : OAI21D0BWP7T port map(A1 => l071_n_91, A2 => l071_n_55, B => l071_n_218, ZN => l071_n_221);
  l071_g12419 : AOI22D0BWP7T port map(A1 => l071_n_205, A2 => l071_n_193, B1 => l071_n_203, B2 => l071_n_178, ZN => l071_n_220);
  l071_g12420 : OAI21D0BWP7T port map(A1 => l071_n_93, A2 => l071_n_64, B => l071_n_217, ZN => l071_n_219);
  l071_g12421 : AOI22D0BWP7T port map(A1 => l071_n_209, A2 => l071_n_151, B1 => l071_n_210, B2 => l071_n_152, ZN => l071_n_225);
  l071_g12422 : OAI32D1BWP7T port map(A1 => l071_n_118, A2 => l071_n_135, A3 => l071_n_198, B1 => l071_n_158, B2 => l071_n_208, ZN => l071_n_223);
  l071_g12423 : AOI22D0BWP7T port map(A1 => l071_n_210, A2 => l071_n_5, B1 => l071_n_209, B2 => l071_n_3, ZN => l071_n_222);
  l071_g12424 : AOI211D1BWP7T port map(A1 => l071_n_128, A2 => l071_n_56, B => l071_n_197, C => l071_n_188, ZN => l071_n_216);
  l071_g12425 : OAI22D0BWP7T port map(A1 => l071_n_200, A2 => l071_n_171, B1 => l071_n_194, B2 => l071_n_181, ZN => l071_n_218);
  l071_g12426 : IOA21D1BWP7T port map(A1 => l071_n_203, A2 => l071_n_167, B => l071_n_211, ZN => l071_n_217);
  l071_g12427 : MOAI22D0BWP7T port map(A1 => l071_n_200, A2 => l071_n_165, B1 => l071_n_203, B2 => l071_n_166, ZN => l071_n_215);
  l071_g12428 : MOAI22D0BWP7T port map(A1 => l071_n_200, A2 => l071_n_168, B1 => l071_n_203, B2 => l071_n_169, ZN => l071_n_214);
  l071_g12429 : MAOI22D0BWP7T port map(A1 => l071_n_201, A2 => l071_n_166, B1 => l071_n_202, B2 => l071_n_165, ZN => l071_n_213);
  l071_g12430 : MOAI22D0BWP7T port map(A1 => l071_n_194, A2 => l071_n_187, B1 => l071_n_201, B2 => l071_n_167, ZN => l071_n_212);
  l071_g12431 : INVD0BWP7T port map(I => l071_n_209, ZN => l071_n_208);
  l071_g12432 : ND2D1BWP7T port map(A1 => l071_n_201, A2 => l071_n_149, ZN => l071_n_211);
  l071_g12433 : NR2D1BWP7T port map(A1 => l071_n_198, A2 => l071_n_113, ZN => l071_n_210);
  l071_g12434 : NR2D1BWP7T port map(A1 => l071_n_198, A2 => l071_n_114, ZN => l071_n_209);
  l071_g12435 : OAI21D0BWP7T port map(A1 => l071_n_131, A2 => l071_n_76, B => l071_n_199, ZN => l071_n_207);
  l071_g12436 : AOI21D0BWP7T port map(A1 => l071_n_143, A2 => l071_n_81, B => l071_n_204, ZN => l071_n_206);
  l071_g12437 : ND4D0BWP7T port map(A1 => l071_n_195, A2 => l071_n_190, A3 => l071_n_2, A4 => l071_n_182, ZN => l071_n_205);
  l071_g12438 : INVD0BWP7T port map(I => l071_n_203, ZN => l071_n_202);
  l071_g12439 : INVD0BWP7T port map(I => l071_n_201, ZN => l071_n_200);
  l071_g12440 : CKND2D1BWP7T port map(A1 => l071_n_193, A2 => l071_n_188, ZN => l071_n_204);
  l071_g12441 : NR2D1BWP7T port map(A1 => l071_n_194, A2 => l071_n_4, ZN => l071_n_203);
  l071_g12442 : NR2D1BWP7T port map(A1 => l071_n_194, A2 => l071_n_185, ZN => l071_n_201);
  l071_g12443 : OA31D1BWP7T port map(A1 => l071_n_120, A2 => l071_n_148, A3 => l071_n_175, B => l071_n_195, Z => l071_n_197);
  l071_g12444 : NR4D0BWP7T port map(A1 => l071_n_194, A2 => l071_n_173, A3 => l071_n_164, A4 => l071_n_43, ZN => l071_n_196);
  l071_g12445 : AOI21D0BWP7T port map(A1 => l071_n_2, A2 => l071_n_182, B => l071_n_194, ZN => l071_n_199);
  l071_g12446 : ND3D0BWP7T port map(A1 => l071_n_193, A2 => l071_n_176, A3 => l071_n_121, ZN => l071_n_198);
  l071_g12447 : INR2XD0BWP7T port map(A1 => l071_n_187, B1 => l071_n_192, ZN => l071_n_195);
  l071_g12448 : INVD1BWP7T port map(I => l071_n_194, ZN => l071_n_193);
  l071_g12449 : OAI221D0BWP7T port map(A1 => l071_n_174, A2 => l071_n_142, B1 => l071_n_29, B2 => l071_n_20, C => l071_n_191, ZN => l071_n_194);
  l071_g12450 : OAI221D0BWP7T port map(A1 => l071_n_185, A2 => l071_n_179, B1 => l071_n_171, B2 => l071_n_4, C => l071_n_181, ZN => l071_n_192);
  l071_g12451 : AOI221D0BWP7T port map(A1 => l071_n_8, A2 => x_enemy1(8), B1 => l071_n_51, B2 => l071_n_17, C => l071_n_186, ZN => l071_n_191);
  l071_g12452 : IAO21D0BWP7T port map(A1 => l071_n_4, A2 => l071_n_183, B => l071_n_189, ZN => l071_n_190);
  l071_g12453 : AOI21D0BWP7T port map(A1 => l071_n_183, A2 => l071_n_171, B => l071_n_185, ZN => l071_n_189);
  l071_g12454 : OAI22D0BWP7T port map(A1 => l071_n_4, A2 => l071_n_168, B1 => l071_n_185, B2 => l071_n_170, ZN => l071_n_188);
  l071_g12455 : IND2D1BWP7T port map(A1 => l071_n_4, B1 => l071_n_149, ZN => l071_n_187);
  l071_g12456 : AO21D0BWP7T port map(A1 => l071_n_20, A2 => l071_n_29, B => l071_n_180, Z => l071_n_186);
  l071_g12458 : NR3D0BWP7T port map(A1 => l071_n_163, A2 => l071_n_91, A3 => l071_n_64, ZN => l071_n_184);
  l071_g12459 : ND2D1BWP7T port map(A1 => l071_n_176, A2 => l071_n_119, ZN => l071_n_185);
  l071_g12461 : MOAI22D0BWP7T port map(A1 => l071_n_51, A2 => l071_n_17, B1 => l071_n_160, B2 => l071_n_142, ZN => l071_n_180);
  l071_g12462 : INR3D0BWP7T port map(A1 => l071_n_168, B1 => l071_n_166, B2 => l071_n_167, ZN => l071_n_183);
  l071_g12463 : ND4D0BWP7T port map(A1 => l071_n_0, A2 => l071_n_155, A3 => l071_n_146, A4 => l071_n_43, ZN => l071_n_182);
  l071_g12464 : IND3D1BWP7T port map(A1 => l071_n_148, B1 => l071_n_120, B2 => l071_n_177, ZN => l071_n_181);
  l071_g12465 : CKND1BWP7T port map(I => l071_n_178, ZN => l071_n_179);
  l071_g12466 : INVD0BWP7T port map(I => l071_n_176, ZN => l071_n_175);
  l071_g12467 : ND2D1BWP7T port map(A1 => l071_n_170, A2 => l071_n_165, ZN => l071_n_178);
  l071_g12468 : AOI211XD0BWP7T port map(A1 => l071_n_46, A2 => l071_n_30, B => l071_n_164, C => l071_n_102, ZN => l071_n_177);
  l071_g12469 : AOI211D1BWP7T port map(A1 => l071_n_46, A2 => l071_n_24, B => l071_n_164, C => l071_n_101, ZN => l071_n_176);
  l071_g12470 : AOI221D0BWP7T port map(A1 => l071_n_107, A2 => l071_n_15, B1 => l071_n_49, B2 => l071_n_105, C => l071_n_159, ZN => l071_n_174);
  l071_g12471 : AOI22D0BWP7T port map(A1 => l071_n_0, A2 => y(4), B1 => l071_n_154, B2 => l071_n_41, ZN => l071_n_173);
  l071_g12472 : INR4D0BWP7T port map(A1 => l071_n_96, B1 => l071_n_94, B2 => l071_n_133, B3 => l071_n_147, ZN => l071_n_172);
  l071_g12473 : INVD0BWP7T port map(I => l071_n_170, ZN => l071_n_169);
  l071_g12474 : ND2D1BWP7T port map(A1 => l071_n_150, A2 => l071_n_113, ZN => l071_n_171);
  l071_g12475 : ND2D1BWP7T port map(A1 => l071_n_152, A2 => l071_n_113, ZN => l071_n_170);
  l071_g12476 : ND2D1BWP7T port map(A1 => l071_n_151, A2 => l071_n_114, ZN => l071_n_168);
  l071_g12477 : INR2D1BWP7T port map(A1 => l071_n_114, B1 => l071_n_158, ZN => l071_n_167);
  l071_g12478 : AN2D1BWP7T port map(A1 => l071_n_5, A2 => l071_n_113, Z => l071_n_166);
  l071_g12479 : ND2D1BWP7T port map(A1 => l071_n_3, A2 => l071_n_114, ZN => l071_n_165);
  l071_g12480 : IND4D0BWP7T port map(A1 => l071_n_71, B1 => l071_n_72, B2 => l071_n_103, B3 => l071_n_116, ZN => l071_n_163);
  l071_g12481 : ND4D0BWP7T port map(A1 => l071_n_129, A2 => l071_n_95, A3 => l071_n_70, A4 => l071_n_60, ZN => l071_n_162);
  l071_g12482 : IND4D0BWP7T port map(A1 => l071_n_76, B1 => l071_n_77, B2 => l071_n_70, B3 => l071_n_124, ZN => l071_n_161);
  l071_g12483 : OAI222D0BWP7T port map(A1 => l071_n_145, A2 => l071_n_138, B1 => l071_n_98, B2 => l071_n_136, C1 => l071_n_105, C2 => l071_n_106, ZN => l071_n_160);
  l071_g12484 : MOAI22D0BWP7T port map(A1 => l071_n_144, A2 => l071_n_137, B1 => l071_n_138, B2 => l071_n_99, ZN => l071_n_159);
  l071_g12485 : ND3D0BWP7T port map(A1 => l071_n_140, A2 => l071_n_146, A3 => l071_n_141, ZN => l071_n_164);
  l071_g12486 : OAI211D1BWP7T port map(A1 => l071_n_13, A2 => l071_n_56, B => l071_n_143, C => l071_n_89, ZN => l071_n_157);
  l071_g12487 : INR3D0BWP7T port map(A1 => l071_n_116, B1 => l071_n_93, B2 => l071_n_125, ZN => l071_n_156);
  l071_g12488 : AOI211D0BWP7T port map(A1 => l071_n_48, A2 => y(5), B => l071_n_123, C => l071_n_109, ZN => l071_n_155);
  l071_g12489 : NR3D0BWP7T port map(A1 => l071_n_134, A2 => l071_n_46, A3 => y(4), ZN => l071_n_154);
  l071_g12490 : AO211D0BWP7T port map(A1 => l071_n_59, A2 => l071_n_11, B => l071_n_147, C => l071_n_86, Z => l071_n_153);
  l071_g12491 : ND3D0BWP7T port map(A1 => l071_n_115, A2 => l071_n_110, A3 => l071_n_45, ZN => l071_n_158);
  l071_g12495 : NR3D0BWP7T port map(A1 => l071_n_117, A2 => l071_n_45, A3 => l071_n_47, ZN => l071_n_152);
  l071_g12496 : NR3D0BWP7T port map(A1 => l071_n_122, A2 => l071_n_115, A3 => l071_n_44, ZN => l071_n_151);
  l071_g12497 : AN4D1BWP7T port map(A1 => l071_n_115, A2 => l071_n_108, A3 => l071_n_1, A4 => l071_n_45, Z => l071_n_150);
  l071_g12498 : INR2D1BWP7T port map(A1 => l071_n_118, B1 => l071_n_135, ZN => l071_n_149);
  l071_g12499 : OR2D1BWP7T port map(A1 => l071_n_134, A2 => l071_n_41, Z => l071_n_148);
  l071_g12500 : ND2D1BWP7T port map(A1 => l071_n_132, A2 => l071_n_95, ZN => l071_n_147);
  l071_g12501 : AOI211XD0BWP7T port map(A1 => l071_n_53, A2 => l071_n_33, B => l071_n_90, C => l071_n_111, ZN => l071_n_146);
  l071_g12502 : CKND1BWP7T port map(I => l071_n_144, ZN => l071_n_145);
  l071_g12503 : AOI22D0BWP7T port map(A1 => l071_n_100, A2 => y(5), B1 => l071_n_83, B2 => y_enemy1(5), ZN => l071_n_141);
  l071_g12504 : NR2D1BWP7T port map(A1 => l071_n_123, A2 => l071_n_109, ZN => l071_n_140);
  l071_g12505 : MAOI222D1BWP7T port map(A => l071_n_88, B => x(2), C => x_enemy1(2), ZN => l071_n_144);
  l071_g12506 : NR3D0BWP7T port map(A1 => l071_n_97, A2 => l071_n_91, A3 => l071_n_69, ZN => l071_n_143);
  l071_g12507 : OAI21D0BWP7T port map(A1 => l071_n_107, A2 => l071_n_14, B => l071_n_106, ZN => l071_n_142);
  l071_g12508 : INVD0BWP7T port map(I => l071_n_136, ZN => l071_n_137);
  l071_g12509 : INVD0BWP7T port map(I => l071_n_132, ZN => l071_n_131);
  l071_g12510 : AOI211XD0BWP7T port map(A1 => l071_n_59, A2 => l071_n_25, B => l071_n_97, C => l071_n_80, ZN => l071_n_130);
  l071_g12511 : OAI21D0BWP7T port map(A1 => l071_n_74, A2 => l071_n_58, B => draw_count5(1), ZN => l071_n_129);
  l071_g12512 : AOI221D0BWP7T port map(A1 => l071_n_58, A2 => l071_n_26, B1 => l071_n_62, B2 => draw_count5(0), C => l071_n_78, ZN => l071_n_128);
  l071_g12513 : AO221D0BWP7T port map(A1 => l071_n_66, A2 => l071_n_64, B1 => l071_n_67, B2 => l071_n_27, C => l071_n_94, Z => l071_n_127);
  l071_g12514 : OA211D0BWP7T port map(A1 => l071_n_25, A2 => l071_n_60, B => l071_n_103, C => l071_n_79, Z => l071_n_126);
  l071_g12515 : OAI211D1BWP7T port map(A1 => l071_n_11, A2 => l071_n_56, B => l071_n_81, C => l071_n_75, ZN => l071_n_125);
  l071_g12516 : AOI21D0BWP7T port map(A1 => l071_n_59, A2 => l071_n_26, B => l071_n_87, ZN => l071_n_124);
  l071_g12517 : AO21D0BWP7T port map(A1 => l071_n_67, A2 => l071_n_66, B => l071_n_94, Z => l071_n_139);
  l071_g12518 : OAI22D0BWP7T port map(A1 => l071_n_68, A2 => l071_n_16, B1 => l071_n_50, B2 => x(2), ZN => l071_n_138);
  l071_g12519 : AOI22D0BWP7T port map(A1 => l071_n_68, A2 => l071_n_16, B1 => l071_n_50, B2 => x(2), ZN => l071_n_136);
  l071_g12520 : ND2D1BWP7T port map(A1 => l071_n_104, A2 => l071_n_42, ZN => l071_n_135);
  l071_g12521 : ND2D1BWP7T port map(A1 => l071_n_104, A2 => l071_n_84, ZN => l071_n_134);
  l071_g12522 : IND2D1BWP7T port map(A1 => l071_n_93, B1 => l071_n_70, ZN => l071_n_133);
  l071_g12523 : INR2XD0BWP7T port map(A1 => l071_n_60, B1 => l071_n_91, ZN => l071_n_132);
  l071_g12528 : OAI22D0BWP7T port map(A1 => l071_n_52, A2 => l071_n_28, B1 => l071_n_48, B2 => y(5), ZN => l071_n_123);
  l071_g12529 : MOAI22D0BWP7T port map(A1 => l071_n_60, A2 => draw_count5(1), B1 => l071_n_74, B2 => l071_n_66, ZN => l071_n_112);
  l071_g12530 : MOAI22D0BWP7T port map(A1 => l071_n_19, A2 => y(9), B1 => l071_n_19, B2 => y(9), ZN => l071_n_111);
  l071_g12531 : MAOI22D0BWP7T port map(A1 => l071_n_84, A2 => l071_n_34, B1 => l071_n_84, B2 => l071_n_34, ZN => l071_n_122);
  l071_g12532 : MAOI22D0BWP7T port map(A1 => l071_n_43, A2 => l071_n_35, B1 => l071_n_43, B2 => l071_n_35, ZN => l071_n_121);
  l071_g12533 : MAOI22D0BWP7T port map(A1 => l071_n_43, A2 => y(3), B1 => l071_n_43, B2 => y(3), ZN => l071_n_120);
  l071_g12534 : MOAI22D0BWP7T port map(A1 => l071_n_43, A2 => l071_n_18, B1 => l071_n_43, B2 => l071_n_18, ZN => l071_n_119);
  l071_g12535 : MAOI22D0BWP7T port map(A1 => l071_n_82, A2 => y(2), B1 => l071_n_82, B2 => y(2), ZN => l071_n_118);
  l071_g12536 : ND2D1BWP7T port map(A1 => l071_n_108, A2 => l071_n_1, ZN => l071_n_110);
  l071_g12537 : MOAI22D0BWP7T port map(A1 => l071_n_42, A2 => y(1), B1 => l071_n_42, B2 => y(1), ZN => l071_n_117);
  l071_g12538 : INR3D0BWP7T port map(A1 => l071_n_79, B1 => l071_n_62, B2 => l071_n_78, ZN => l071_n_116);
  l071_g12539 : MOAI22D0BWP7T port map(A1 => l071_n_47, A2 => y(0), B1 => l071_n_47, B2 => y(0), ZN => l071_n_115);
  l071_g12540 : MAOI22D0BWP7T port map(A1 => l071_n_41, A2 => l071_n_21, B1 => l071_n_41, B2 => l071_n_21, ZN => l071_n_114);
  l071_g12541 : MOAI22D0BWP7T port map(A1 => l071_n_41, A2 => l071_n_23, B1 => l071_n_41, B2 => l071_n_23, ZN => l071_n_113);
  l071_g12542 : NR2XD0BWP7T port map(A1 => l071_n_46, A2 => l071_n_30, ZN => l071_n_102);
  l071_g12543 : NR2XD0BWP7T port map(A1 => l071_n_46, A2 => l071_n_24, ZN => l071_n_101);
  l071_g12545 : CKAN2D1BWP7T port map(A1 => l071_n_52, A2 => l071_n_28, Z => l071_n_109);
  l071_g12546 : ND2D1BWP7T port map(A1 => l071_n_42, A2 => l071_n_31, ZN => l071_n_108);
  l071_g12547 : NR2XD0BWP7T port map(A1 => l071_n_83, A2 => y_enemy1(5), ZN => l071_n_100);
  l071_g12548 : CKAN2D1BWP7T port map(A1 => l071_n_49, A2 => l071_n_38, Z => l071_n_107);
  l071_g12550 : OR2D1BWP7T port map(A1 => l071_n_49, A2 => l071_n_15, Z => l071_n_106);
  l071_g12551 : NR2XD0BWP7T port map(A1 => l071_n_68, A2 => l071_n_16, ZN => l071_n_98);
  l071_g12552 : AN2D0BWP7T port map(A1 => l071_n_14, A2 => l071_n_38, Z => l071_n_105);
  l071_g12553 : INR2D1BWP7T port map(A1 => l071_n_47, B1 => l071_n_45, ZN => l071_n_104);
  l071_g12554 : NR2XD0BWP7T port map(A1 => l071_n_73, A2 => l071_n_80, ZN => l071_n_103);
  l071_g12555 : NR2D1BWP7T port map(A1 => l071_n_53, A2 => l071_n_33, ZN => l071_n_90);
  l071_g12556 : AOI22D0BWP7T port map(A1 => l071_n_59, A2 => l071_n_12, B1 => l071_n_62, B2 => l071_n_25, ZN => l071_n_89);
  l071_g12557 : AOI22D0BWP7T port map(A1 => l071_n_54, A2 => x(0), B1 => x(1), B2 => l071_n_9, ZN => l071_n_88);
  l071_g12558 : AOI21D0BWP7T port map(A1 => l071_n_57, A2 => l071_n_60, B => draw_count5(1), ZN => l071_n_87);
  l071_g12559 : OA21D0BWP7T port map(A1 => l071_n_58, A2 => l071_n_55, B => l071_n_25, Z => l071_n_86);
  l071_g12560 : AOI21D0BWP7T port map(A1 => l071_n_58, A2 => l071_n_25, B => l071_n_63, ZN => l071_n_85);
  l071_g12561 : OAI21D0BWP7T port map(A1 => l071_n_56, A2 => draw_count5(1), B => l071_n_75, ZN => l071_n_97);
  l071_g12562 : AOI21D0BWP7T port map(A1 => l071_n_62, A2 => l071_n_11, B => l071_n_59, ZN => l071_n_96);
  l071_g12563 : OAI21D0BWP7T port map(A1 => l071_n_63, A2 => l071_n_55, B => l071_n_12, ZN => l071_n_95);
  l071_g12564 : MOAI22D0BWP7T port map(A1 => l071_n_65, A2 => l071_n_26, B1 => l071_n_67, B2 => l071_n_12, ZN => l071_n_94);
  l071_g12565 : AO21D0BWP7T port map(A1 => l071_n_64, A2 => l071_n_26, B => l071_n_73, Z => l071_n_93);
  l071_g12566 : IOA21D1BWP7T port map(A1 => l071_n_58, A2 => l071_n_11, B => l071_n_77, ZN => l071_n_92);
  l071_g12567 : OAI22D0BWP7T port map(A1 => l071_n_57, A2 => l071_n_11, B1 => l071_n_60, B2 => l071_n_26, ZN => l071_n_91);
  l071_g12568 : INVD1BWP7T port map(I => l071_n_42, ZN => l071_n_84);
  l071_g12570 : INVD0BWP7T port map(I => l071_n_48, ZN => l071_n_83);
  l071_g12571 : INVD0BWP7T port map(I => l071_n_41, ZN => l071_n_82);
  l071_g12572 : ND2D1BWP7T port map(A1 => l071_n_59, A2 => draw_count5(1), ZN => l071_n_81);
  l071_g12573 : NR2D1BWP7T port map(A1 => l071_n_65, A2 => draw_count5(1), ZN => l071_n_80);
  l071_g12574 : IND2D0BWP7T port map(A1 => l071_n_13, B1 => l071_n_63, ZN => l071_n_79);
  l071_g12575 : INR2D1BWP7T port map(A1 => l071_n_59, B1 => draw_count5(1), ZN => l071_n_78);
  l071_g12576 : CKND2D0BWP7T port map(A1 => l071_n_63, A2 => l071_n_12, ZN => l071_n_77);
  l071_g12577 : NR2D0BWP7T port map(A1 => l071_n_56, A2 => l071_n_6, ZN => l071_n_76);
  l071_g12578 : NR2D0BWP7T port map(A1 => l071_n_60, A2 => l071_n_13, ZN => l071_n_69);
  l071_g12579 : CKND2D1BWP7T port map(A1 => l071_n_58, A2 => l071_n_66, ZN => l071_n_75);
  l071_g12580 : IND2D1BWP7T port map(A1 => l071_n_59, B1 => l071_n_61, ZN => l071_n_74);
  l071_g12581 : AN2D0BWP7T port map(A1 => l071_n_63, A2 => l071_n_25, Z => l071_n_73);
  l071_g12582 : ND2D1BWP7T port map(A1 => l071_n_55, A2 => l071_n_11, ZN => l071_n_72);
  l071_g12583 : INR2D1BWP7T port map(A1 => l071_n_27, B1 => l071_n_57, ZN => l071_n_71);
  l071_g12584 : ND2D1BWP7T port map(A1 => l071_n_63, A2 => l071_n_66, ZN => l071_n_70);
  l071_g12585 : INVD1BWP7T port map(I => l071_n_65, ZN => l071_n_64);
  l071_g12586 : INVD1BWP7T port map(I => l071_n_62, ZN => l071_n_61);
  l071_g12587 : INVD0BWP7T port map(I => l071_n_58, ZN => l071_n_57);
  l071_g12588 : INVD1BWP7T port map(I => l071_n_56, ZN => l071_n_55);
  l071_g12589 : IAO21D0BWP7T port map(A1 => x(1), A2 => l071_n_9, B => x_enemy1(0), ZN => l071_n_54);
  l071_g12590 : AO21D0BWP7T port map(A1 => x(4), A2 => l071_n_10, B => l071_n_14, Z => l071_n_68);
  l071_g12591 : INR2D1BWP7T port map(A1 => draw_count5(3), B1 => l071_n_32, ZN => l071_n_67);
  l071_g12592 : IND2D1BWP7T port map(A1 => l071_n_27, B1 => l071_n_13, ZN => l071_n_66);
  l071_g12593 : ND2D1BWP7T port map(A1 => l071_n_39, A2 => draw_count5(3), ZN => l071_n_65);
  l071_g12594 : NR2D1BWP7T port map(A1 => l071_n_32, A2 => draw_count5(3), ZN => l071_n_63);
  l071_g12595 : INR2D1BWP7T port map(A1 => l071_n_22, B1 => draw_count5(3), ZN => l071_n_62);
  l071_g12596 : ND2D1BWP7T port map(A1 => l071_n_36, A2 => draw_count5(3), ZN => l071_n_60);
  l071_g12597 : NR2D1BWP7T port map(A1 => l071_n_37, A2 => draw_count5(3), ZN => l071_n_59);
  l071_g12598 : NR2D1BWP7T port map(A1 => l071_n_40, A2 => draw_count5(3), ZN => l071_n_58);
  l071_g12599 : ND2D1BWP7T port map(A1 => l071_n_22, A2 => draw_count5(3), ZN => l071_n_56);
  l071_g12601 : INVD0BWP7T port map(I => l071_n_45, ZN => l071_n_44);
  l071_g12602 : MOAI22D0BWP7T port map(A1 => y(8), A2 => y_enemy1(8), B1 => y(8), B2 => y_enemy1(8), ZN => l071_n_53);
  l071_g12603 : MAOI22D0BWP7T port map(A1 => y(7), A2 => y_enemy1(7), B1 => y(7), B2 => y_enemy1(7), ZN => l071_n_52);
  l071_g12604 : MOAI22D0BWP7T port map(A1 => x(7), A2 => x_enemy1(7), B1 => x(7), B2 => x_enemy1(7), ZN => l071_n_51);
  l071_g12605 : MAOI22D0BWP7T port map(A1 => x(3), A2 => x_enemy1(3), B1 => x(3), B2 => x_enemy1(3), ZN => l071_n_50);
  l071_g12606 : MAOI22D0BWP7T port map(A1 => x(6), A2 => x_enemy1(6), B1 => x(6), B2 => x_enemy1(6), ZN => l071_n_49);
  l071_g12607 : OAI21D0BWP7T port map(A1 => l071_n_7, A2 => y_enemy1(6), B => l071_n_28, ZN => l071_n_48);
  l071_g12608 : MOAI22D0BWP7T port map(A1 => y(1), A2 => y_enemy1(1), B1 => y(1), B2 => y_enemy1(1), ZN => l071_n_47);
  l071_g12609 : MAOI22D0BWP7T port map(A1 => y(5), A2 => y_enemy1(5), B1 => y(5), B2 => y_enemy1(5), ZN => l071_n_46);
  l071_g12610 : MAOI22D0BWP7T port map(A1 => y(0), A2 => y_enemy1(0), B1 => y(0), B2 => y_enemy1(0), ZN => l071_n_45);
  l071_g12611 : MOAI22D0BWP7T port map(A1 => y(4), A2 => y_enemy1(4), B1 => y(4), B2 => y_enemy1(4), ZN => l071_n_43);
  l071_g12612 : MAOI22D0BWP7T port map(A1 => y(2), A2 => y_enemy1(2), B1 => y(2), B2 => y_enemy1(2), ZN => l071_n_42);
  l071_g12613 : MOAI22D0BWP7T port map(A1 => y(3), A2 => y_enemy1(3), B1 => y(3), B2 => y_enemy1(3), ZN => l071_n_41);
  l071_g12614 : INVD0BWP7T port map(I => l071_n_39, ZN => l071_n_40);
  l071_g12615 : CKND1BWP7T port map(I => l071_n_36, ZN => l071_n_37);
  l071_g12616 : INVD1BWP7T port map(I => l071_n_26, ZN => l071_n_25);
  l071_g12617 : INR2D1BWP7T port map(A1 => draw_count5(4), B1 => draw_count5(2), ZN => l071_n_39);
  l071_g12618 : IND2D0BWP7T port map(A1 => x_enemy1(5), B1 => x(5), ZN => l071_n_38);
  l071_g12619 : INR2D1BWP7T port map(A1 => draw_count5(2), B1 => draw_count5(4), ZN => l071_n_36);
  l071_g12620 : IND2D0BWP7T port map(A1 => y_enemy1(3), B1 => y(3), ZN => l071_n_35);
  l071_g12621 : IND2D1BWP7T port map(A1 => y_enemy1(1), B1 => y(1), ZN => l071_n_34);
  l071_g12622 : INR2XD0BWP7T port map(A1 => y_enemy1(7), B1 => y(7), ZN => l071_n_33);
  l071_g12623 : ND2D1BWP7T port map(A1 => draw_count5(2), A2 => draw_count5(4), ZN => l071_n_32);
  l071_g12624 : IND2D1BWP7T port map(A1 => y(1), B1 => y_enemy1(1), ZN => l071_n_31);
  l071_g12625 : IND2D0BWP7T port map(A1 => y_enemy1(4), B1 => y(4), ZN => l071_n_30);
  l071_g12626 : IND2D1BWP7T port map(A1 => x(7), B1 => x_enemy1(7), ZN => l071_n_29);
  l071_g12627 : ND2D1BWP7T port map(A1 => l071_n_7, A2 => y_enemy1(6), ZN => l071_n_28);
  l071_g12628 : INR2D1BWP7T port map(A1 => draw_count5(0), B1 => draw_count5(1), ZN => l071_n_27);
  l071_g12629 : CKND2D1BWP7T port map(A1 => draw_count5(1), A2 => draw_count5(0), ZN => l071_n_26);
  l071_g12630 : INVD1BWP7T port map(I => l071_n_12, ZN => l071_n_11);
  l071_g12631 : INR2XD0BWP7T port map(A1 => y_enemy1(4), B1 => y(4), ZN => l071_n_24);
  l071_g12632 : IND2D1BWP7T port map(A1 => y(2), B1 => y_enemy1(2), ZN => l071_n_23);
  l071_g12633 : NR2D0BWP7T port map(A1 => draw_count5(2), A2 => draw_count5(4), ZN => l071_n_22);
  l071_g12634 : IND2D1BWP7T port map(A1 => y_enemy1(2), B1 => y(2), ZN => l071_n_21);
  l071_g12635 : NR2D1BWP7T port map(A1 => l071_n_8, A2 => x_enemy1(8), ZN => l071_n_20);
  l071_g12636 : IND2D1BWP7T port map(A1 => y(8), B1 => y_enemy1(8), ZN => l071_n_19);
  l071_g12637 : IND2D1BWP7T port map(A1 => y(3), B1 => y_enemy1(3), ZN => l071_n_18);
  l071_g12638 : IND2D1BWP7T port map(A1 => x_enemy1(6), B1 => x(6), ZN => l071_n_17);
  l071_g12639 : IND2D1BWP7T port map(A1 => x(3), B1 => x_enemy1(3), ZN => l071_n_16);
  l071_g12640 : INR2XD0BWP7T port map(A1 => x_enemy1(5), B1 => x(5), ZN => l071_n_15);
  l071_g12641 : NR2D0BWP7T port map(A1 => x(4), A2 => l071_n_10, ZN => l071_n_14);
  l071_g12642 : IND2D1BWP7T port map(A1 => draw_count5(0), B1 => draw_count5(1), ZN => l071_n_13);
  l071_g12643 : NR2D0BWP7T port map(A1 => draw_count5(1), A2 => draw_count5(0), ZN => l071_n_12);
  l071_g12644 : CKND1BWP7T port map(I => x_enemy1(4), ZN => l071_n_10);
  l071_g12645 : INVD0BWP7T port map(I => x_enemy1(1), ZN => l071_n_9);
  l071_g12646 : CKND1BWP7T port map(I => x(8), ZN => l071_n_8);
  l071_g12647 : CKND1BWP7T port map(I => y(6), ZN => l071_n_7);
  l071_g12648 : INVD0BWP7T port map(I => draw_count5(1), ZN => l071_n_6);
  l071_g2 : INR3D0BWP7T port map(A1 => l071_n_122, B1 => l071_n_115, B2 => l071_n_44, ZN => l071_n_5);
  l071_g12649 : IND2D1BWP7T port map(A1 => l071_n_119, B1 => l071_n_177, ZN => l071_n_4);
  l071_g12650 : INR3D0BWP7T port map(A1 => l071_n_117, B1 => l071_n_45, B2 => l071_n_47, ZN => l071_n_3);
  l071_g12651 : IIND4D0BWP7T port map(A1 => l071_n_121, A2 => l071_n_113, B1 => l071_n_150, B2 => l071_n_177, ZN => l071_n_2);
  l071_g12652 : IND2D1BWP7T port map(A1 => l071_n_31, B1 => l071_n_84, ZN => l071_n_1);
  l071_g12653 : INR3D0BWP7T port map(A1 => l071_n_46, B1 => l071_n_134, B2 => l071_n_82, ZN => l071_n_0);
  l071_g12654 : INVD0BWP7T port map(I => l071_n_68, ZN => l071_n_99);
  l053_g2484 : OA21D0BWP7T port map(A1 => l053_n_82, A2 => l053_n_39, B => enable3, Z => r3);
  l053_g2485 : AO31D1BWP7T port map(A1 => l053_n_79, A2 => l053_n_77, A3 => draw_count3(0), B => b3, Z => g3);
  l053_g2486 : AO31D1BWP7T port map(A1 => l053_n_79, A2 => l053_n_77, A3 => l053_n_15, B => l053_n_83, Z => b3);
  l053_g2487 : OA21D0BWP7T port map(A1 => l053_n_80, A2 => l053_n_78, B => l053_n_39, Z => l053_n_83);
  l053_g2488 : OAI22D0BWP7T port map(A1 => l053_n_80, A2 => l053_n_73, B1 => l053_n_2, B2 => draw_count3(2), ZN => l053_n_82);
  l053_g2489 : OR2D1BWP7T port map(A1 => l053_n_77, A2 => l053_n_78, Z => enable3);
  l053_g2490 : INVD0BWP7T port map(I => l053_n_80, ZN => l053_n_79);
  l053_g2491 : NR2D1BWP7T port map(A1 => l053_n_76, A2 => l053_n_74, ZN => l053_n_80);
  l053_g2492 : INR2D1BWP7T port map(A1 => l053_n_73, B1 => l053_n_76, ZN => l053_n_78);
  l053_g2493 : AOI21D0BWP7T port map(A1 => l053_n_74, A2 => l053_n_0, B => l053_n_76, ZN => l053_n_77);
  l053_g2494 : OAI221D0BWP7T port map(A1 => l053_n_31, A2 => l053_n_9, B1 => l053_n_10, B2 => l053_n_33, C => l053_n_75, ZN => l053_n_76);
  l053_g2495 : NR4D0BWP7T port map(A1 => l053_n_71, A2 => l053_n_67, A3 => l053_n_60, A4 => l053_n_53, ZN => l053_n_75);
  l053_g2497 : ND4D0BWP7T port map(A1 => l053_n_72, A2 => l053_n_57, A3 => l053_n_35, A4 => l053_n_29, ZN => l053_n_74);
  l053_g2498 : NR4D0BWP7T port map(A1 => l053_n_70, A2 => l053_n_35, A3 => l053_n_36, A4 => l053_n_26, ZN => l053_n_73);
  l053_g2499 : AOI211XD0BWP7T port map(A1 => l053_n_30, A2 => l053_n_16, B => l053_n_69, C => l053_n_63, ZN => l053_n_72);
  l053_g2500 : OAI211D1BWP7T port map(A1 => l053_n_14, A2 => l053_n_25, B => l053_n_68, C => l053_n_51, ZN => l053_n_71);
  l053_g2501 : ND4D0BWP7T port map(A1 => l053_n_65, A2 => l053_n_61, A3 => l053_n_37, A4 => l053_n_29, ZN => l053_n_70);
  l053_g2502 : OAI211D1BWP7T port map(A1 => l053_n_16, A2 => l053_n_30, B => l053_n_66, C => l053_n_56, ZN => l053_n_69);
  l053_g2503 : MAOI222D1BWP7T port map(A => l053_n_64, B => l053_n_34, C => l053_n_5, ZN => l053_n_68);
  l053_g2504 : AOI22D0BWP7T port map(A1 => l053_n_62, A2 => l053_n_52, B1 => l053_n_34, B2 => l053_n_18, ZN => l053_n_67);
  l053_g2505 : AN3D1BWP7T port map(A1 => l053_n_55, A2 => l053_n_50, A3 => l053_n_61, Z => l053_n_66);
  l053_g2506 : NR3D0BWP7T port map(A1 => l053_n_63, A2 => l053_n_54, A3 => l053_n_30, ZN => l053_n_65);
  l053_g2507 : MAOI222D1BWP7T port map(A => l053_n_48, B => l053_n_28, C => x(2), ZN => l053_n_64);
  l053_g2508 : OAI211D1BWP7T port map(A1 => l053_n_17, A2 => l053_n_32, B => l053_n_47, C => l053_n_59, ZN => l053_n_63);
  l053_g2509 : AO211D0BWP7T port map(A1 => l053_n_28, A2 => l053_n_19, B => l053_n_46, C => l053_n_42, Z => l053_n_62);
  l053_g2510 : MOAI22D0BWP7T port map(A1 => x(8), A2 => l053_n_1, B1 => l053_n_31, B2 => l053_n_9, ZN => l053_n_60);
  l053_g2511 : MAOI22D0BWP7T port map(A1 => l053_n_20, A2 => y(9), B1 => l053_n_20, B2 => y(9), ZN => l053_n_59);
  l053_g2512 : MAOI22D0BWP7T port map(A1 => l053_n_26, A2 => l053_n_13, B1 => l053_n_26, B2 => l053_n_13, ZN => l053_n_58);
  l053_g2513 : MAOI22D0BWP7T port map(A1 => l053_n_26, A2 => y(1), B1 => l053_n_26, B2 => y(1), ZN => l053_n_57);
  l053_g2514 : MAOI22D0BWP7T port map(A1 => l053_n_37, A2 => l053_n_11, B1 => l053_n_37, B2 => l053_n_11, ZN => l053_n_56);
  l053_g2515 : MOAI22D0BWP7T port map(A1 => l053_n_38, A2 => l053_n_12, B1 => l053_n_38, B2 => l053_n_12, ZN => l053_n_61);
  l053_g2516 : MAOI22D0BWP7T port map(A1 => l053_n_45, A2 => l053_n_44, B1 => l053_n_36, B2 => l053_n_22, ZN => l053_n_55);
  l053_g2517 : MOAI22D0BWP7T port map(A1 => l053_n_45, A2 => y(5), B1 => l053_n_45, B2 => y(5), ZN => l053_n_54);
  l053_g2518 : MOAI22D0BWP7T port map(A1 => l053_n_40, A2 => l053_n_24, B1 => l053_n_14, B2 => l053_n_25, ZN => l053_n_53);
  l053_g2519 : OA22D0BWP7T port map(A1 => l053_n_34, A2 => l053_n_18, B1 => l053_n_19, B2 => l053_n_28, Z => l053_n_52);
  l053_g2520 : AOI22D0BWP7T port map(A1 => l053_n_40, A2 => l053_n_24, B1 => l053_n_33, B2 => l053_n_10, ZN => l053_n_51);
  l053_g2521 : AOI22D0BWP7T port map(A1 => l053_n_36, A2 => l053_n_22, B1 => l053_n_27, B2 => l053_n_7, ZN => l053_n_50);
  l053_g2522 : MAOI22D0BWP7T port map(A1 => l053_n_35, A2 => y(0), B1 => l053_n_35, B2 => y(0), ZN => l053_n_49);
  l053_g2523 : OR2D1BWP7T port map(A1 => l053_n_43, A2 => l053_n_6, Z => l053_n_48);
  l053_g2524 : ND2D1BWP7T port map(A1 => l053_n_32, A2 => l053_n_17, ZN => l053_n_47);
  l053_g2525 : OA21D0BWP7T port map(A1 => l053_n_41, A2 => l053_n_6, B => l053_n_23, Z => l053_n_46);
  l053_g2526 : INVD0BWP7T port map(I => l053_n_27, ZN => l053_n_45);
  l053_g2527 : INVD0BWP7T port map(I => l053_n_7, ZN => l053_n_44);
  l053_g2528 : AOI21D0BWP7T port map(A1 => l053_n_21, A2 => l053_n_23, B => l053_n_41, ZN => l053_n_43);
  l053_g2529 : OA21D0BWP7T port map(A1 => l053_n_8, A2 => l053_n_6, B => l053_n_21, Z => l053_n_42);
  l053_g2530 : AO21D0BWP7T port map(A1 => l053_n_4, A2 => x_bullet3(1), B => l053_n_8, Z => l053_n_41);
  l053_g2531 : MAOI22D0BWP7T port map(A1 => x(6), A2 => x_bullet3(6), B1 => x(6), B2 => x_bullet3(6), ZN => l053_n_40);
  l053_g2532 : OA21D0BWP7T port map(A1 => l053_n_2, A2 => draw_count3(1), B => l053_n_15, Z => l053_n_39);
  l053_g2533 : MOAI22D0BWP7T port map(A1 => y(7), A2 => y_bullet3(7), B1 => y(7), B2 => y_bullet3(7), ZN => l053_n_38);
  l053_g2534 : OAI21D0BWP7T port map(A1 => y(5), A2 => l053_n_3, B => l053_n_7, ZN => l053_n_37);
  l053_g2535 : MAOI22D0BWP7T port map(A1 => y(4), A2 => y_bullet3(4), B1 => y(4), B2 => y_bullet3(4), ZN => l053_n_36);
  l053_g2536 : MAOI22D0BWP7T port map(A1 => y(1), A2 => y_bullet3(1), B1 => y(1), B2 => y_bullet3(1), ZN => l053_n_35);
  l053_g2537 : MOAI22D0BWP7T port map(A1 => x(4), A2 => x_bullet3(4), B1 => x(4), B2 => x_bullet3(4), ZN => l053_n_34);
  l053_g2539 : MOAI22D0BWP7T port map(A1 => x(5), A2 => x_bullet3(5), B1 => x(5), B2 => x_bullet3(5), ZN => l053_n_33);
  l053_g2540 : MOAI22D0BWP7T port map(A1 => y(8), A2 => y_bullet3(8), B1 => y(8), B2 => y_bullet3(8), ZN => l053_n_32);
  l053_g2541 : MOAI22D0BWP7T port map(A1 => x(7), A2 => x_bullet3(7), B1 => x(7), B2 => x_bullet3(7), ZN => l053_n_31);
  l053_g2542 : MAOI22D0BWP7T port map(A1 => y(3), A2 => y_bullet3(3), B1 => y(3), B2 => y_bullet3(3), ZN => l053_n_30);
  l053_g2543 : MOAI22D0BWP7T port map(A1 => y(0), A2 => y_bullet3(0), B1 => y(0), B2 => y_bullet3(0), ZN => l053_n_29);
  l053_g2544 : MAOI22D0BWP7T port map(A1 => x(3), A2 => x_bullet3(3), B1 => x(3), B2 => x_bullet3(3), ZN => l053_n_28);
  l053_g2545 : MOAI22D0BWP7T port map(A1 => y(6), A2 => y_bullet3(6), B1 => y(6), B2 => y_bullet3(6), ZN => l053_n_27);
  l053_g2546 : MAOI22D0BWP7T port map(A1 => y(2), A2 => y_bullet3(2), B1 => y(2), B2 => y_bullet3(2), ZN => l053_n_26);
  l053_g2547 : IND2D1BWP7T port map(A1 => x(7), B1 => x_bullet3(7), ZN => l053_n_25);
  l053_g2548 : INR2D0BWP7T port map(A1 => x_bullet3(5), B1 => x(5), ZN => l053_n_24);
  l053_g2549 : IND2D0BWP7T port map(A1 => x_bullet3(0), B1 => x(0), ZN => l053_n_23);
  l053_g2550 : IND2D1BWP7T port map(A1 => y(3), B1 => y_bullet3(3), ZN => l053_n_22);
  l053_g2551 : IND2D0BWP7T port map(A1 => x_bullet3(1), B1 => x(1), ZN => l053_n_21);
  l053_g2552 : IND2D1BWP7T port map(A1 => y(8), B1 => y_bullet3(8), ZN => l053_n_20);
  l053_g2553 : INR2D0BWP7T port map(A1 => x_bullet3(2), B1 => x(2), ZN => l053_n_19);
  l053_g2554 : IND2D0BWP7T port map(A1 => x_bullet3(3), B1 => x(3), ZN => l053_n_18);
  l053_g2555 : INR2XD0BWP7T port map(A1 => y_bullet3(7), B1 => y(7), ZN => l053_n_17);
  l053_g2556 : IND2D1BWP7T port map(A1 => y(2), B1 => y_bullet3(2), ZN => l053_n_16);
  l053_g2557 : OR2D1BWP7T port map(A1 => draw_count3(1), A2 => draw_count3(2), Z => l053_n_15);
  l053_g2558 : AN2D1BWP7T port map(A1 => x(8), A2 => l053_n_1, Z => l053_n_14);
  l053_g2559 : INR2D0BWP7T port map(A1 => x_bullet3(3), B1 => x(3), ZN => l053_n_5);
  l053_g2560 : IND2D1BWP7T port map(A1 => y(1), B1 => y_bullet3(1), ZN => l053_n_13);
  l053_g2561 : IND2D1BWP7T port map(A1 => y(6), B1 => y_bullet3(6), ZN => l053_n_12);
  l053_g2562 : INR2XD0BWP7T port map(A1 => y_bullet3(4), B1 => y(4), ZN => l053_n_11);
  l053_g2563 : INR2D0BWP7T port map(A1 => x_bullet3(4), B1 => x(4), ZN => l053_n_10);
  l053_g2564 : IND2D0BWP7T port map(A1 => x_bullet3(6), B1 => x(6), ZN => l053_n_9);
  l053_g2565 : AN2D0BWP7T port map(A1 => x(2), A2 => x_bullet3(2), Z => l053_n_8);
  l053_g2566 : ND2D1BWP7T port map(A1 => y(5), A2 => l053_n_3, ZN => l053_n_7);
  l053_g2567 : NR2D0BWP7T port map(A1 => x(2), A2 => x_bullet3(2), ZN => l053_n_6);
  l053_g2568 : INVD0BWP7T port map(I => x(1), ZN => l053_n_4);
  l053_g2569 : INVD1BWP7T port map(I => y_bullet3(5), ZN => l053_n_3);
  l053_g2570 : INVD0BWP7T port map(I => draw_count3(0), ZN => l053_n_2);
  l053_g2571 : INVD0BWP7T port map(I => x_bullet3(8), ZN => l053_n_1);
  l053_g2 : IND4D0BWP7T port map(A1 => l053_n_29, B1 => l053_n_72, B2 => l053_n_49, B3 => l053_n_58, ZN => l053_n_0);
  l072_g12419 : OAI221D0BWP7T port map(A1 => l072_n_222, A2 => l072_n_184, B1 => l072_n_156, B2 => l072_n_225, C => l072_n_246, ZN => r6);
  l072_g12420 : NR4D0BWP7T port map(A1 => l072_n_245, A2 => l072_n_235, A3 => l072_n_229, A4 => l072_n_206, ZN => l072_n_246);
  l072_g12421 : IND4D0BWP7T port map(A1 => l072_n_233, B1 => l072_n_228, B2 => l072_n_234, B3 => l072_n_242, ZN => l072_n_245);
  l072_g12422 : AO211D0BWP7T port map(A1 => l072_n_218, A2 => l072_n_92, B => l072_n_243, C => l072_n_241, Z => g6);
  l072_g12423 : OAI211D1BWP7T port map(A1 => l072_n_126, A2 => l072_n_222, B => l072_n_239, C => l072_n_231, ZN => l072_n_243);
  l072_g12424 : MAOI22D0BWP7T port map(A1 => l072_n_215, A2 => l072_n_162, B1 => l072_n_236, B2 => l072_n_194, ZN => l072_n_242);
  l072_g12425 : AO221D0BWP7T port map(A1 => l072_n_215, A2 => l072_n_139, B1 => l072_n_212, B2 => l072_n_127, C => l072_n_237, Z => l072_n_241);
  l072_g12426 : OAI32D1BWP7T port map(A1 => l072_n_25, A2 => l072_n_61, A3 => l072_n_222, B1 => l072_n_96, B2 => l072_n_224, ZN => b6);
  l072_g12427 : AOI211XD0BWP7T port map(A1 => l072_n_199, A2 => l072_n_71, B => l072_n_232, C => l072_n_226, ZN => l072_n_239);
  l072_g12428 : ND3D0BWP7T port map(A1 => l072_n_220, A2 => l072_n_211, A3 => l072_n_198, ZN => enable6);
  l072_g12429 : OAI211D1BWP7T port map(A1 => l072_n_85, A2 => l072_n_204, B => l072_n_219, C => l072_n_227, ZN => l072_n_237);
  l072_g12430 : ND4D0BWP7T port map(A1 => l072_n_216, A2 => l072_n_187, A3 => l072_n_181, A4 => l072_n_165, ZN => l072_n_236);
  l072_g12431 : OAI211D1BWP7T port map(A1 => l072_n_172, A2 => l072_n_224, B => l072_n_221, C => l072_n_207, ZN => l072_n_235);
  l072_g12432 : AOI22D0BWP7T port map(A1 => l072_n_212, A2 => l072_n_157, B1 => l072_n_217, B2 => l072_n_161, ZN => l072_n_234);
  l072_g12433 : AOI31D0BWP7T port map(A1 => l072_n_130, A2 => l072_n_132, A3 => l072_n_61, B => l072_n_230, ZN => l072_n_233);
  l072_g12434 : AOI21D0BWP7T port map(A1 => l072_n_132, A2 => l072_n_72, B => l072_n_225, ZN => l072_n_232);
  l072_g12435 : OAI21D0BWP7T port map(A1 => l072_n_133, A2 => l072_n_92, B => l072_n_223, ZN => l072_n_231);
  l072_g12436 : AOI21D0BWP7T port map(A1 => l072_n_210, A2 => l072_n_150, B => l072_n_196, ZN => l072_n_230);
  l072_g12437 : IAO21D0BWP7T port map(A1 => l072_n_153, A2 => l072_n_71, B => l072_n_213, ZN => l072_n_229);
  l072_g12438 : OAI31D0BWP7T port map(A1 => l072_n_76, A2 => l072_n_92, A3 => l072_n_112, B => l072_n_214, ZN => l072_n_228);
  l072_g12439 : OAI21D0BWP7T port map(A1 => l072_n_133, A2 => l072_n_139, B => l072_n_214, ZN => l072_n_227);
  l072_g12440 : AOI21D0BWP7T port map(A1 => l072_n_102, A2 => l072_n_70, B => l072_n_213, ZN => l072_n_226);
  l072_g12441 : INVD0BWP7T port map(I => l072_n_223, ZN => l072_n_224);
  l072_g12442 : OAI21D0BWP7T port map(A1 => l072_n_91, A2 => l072_n_55, B => l072_n_218, ZN => l072_n_221);
  l072_g12443 : AOI22D0BWP7T port map(A1 => l072_n_205, A2 => l072_n_193, B1 => l072_n_203, B2 => l072_n_178, ZN => l072_n_220);
  l072_g12444 : OAI21D0BWP7T port map(A1 => l072_n_93, A2 => l072_n_64, B => l072_n_217, ZN => l072_n_219);
  l072_g12445 : AOI22D0BWP7T port map(A1 => l072_n_209, A2 => l072_n_151, B1 => l072_n_210, B2 => l072_n_3, ZN => l072_n_225);
  l072_g12446 : OAI32D1BWP7T port map(A1 => l072_n_118, A2 => l072_n_135, A3 => l072_n_198, B1 => l072_n_158, B2 => l072_n_208, ZN => l072_n_223);
  l072_g12447 : AOI22D0BWP7T port map(A1 => l072_n_210, A2 => l072_n_5, B1 => l072_n_209, B2 => l072_n_152, ZN => l072_n_222);
  l072_g12448 : AOI211D1BWP7T port map(A1 => l072_n_128, A2 => l072_n_56, B => l072_n_197, C => l072_n_188, ZN => l072_n_216);
  l072_g12449 : OAI22D0BWP7T port map(A1 => l072_n_200, A2 => l072_n_171, B1 => l072_n_194, B2 => l072_n_181, ZN => l072_n_218);
  l072_g12450 : IOA21D1BWP7T port map(A1 => l072_n_203, A2 => l072_n_167, B => l072_n_211, ZN => l072_n_217);
  l072_g12451 : MOAI22D0BWP7T port map(A1 => l072_n_200, A2 => l072_n_165, B1 => l072_n_203, B2 => l072_n_166, ZN => l072_n_215);
  l072_g12452 : MOAI22D0BWP7T port map(A1 => l072_n_200, A2 => l072_n_168, B1 => l072_n_203, B2 => l072_n_169, ZN => l072_n_214);
  l072_g12453 : MAOI22D0BWP7T port map(A1 => l072_n_201, A2 => l072_n_166, B1 => l072_n_202, B2 => l072_n_165, ZN => l072_n_213);
  l072_g12454 : MOAI22D0BWP7T port map(A1 => l072_n_194, A2 => l072_n_187, B1 => l072_n_201, B2 => l072_n_167, ZN => l072_n_212);
  l072_g12455 : INVD0BWP7T port map(I => l072_n_209, ZN => l072_n_208);
  l072_g12456 : ND2D1BWP7T port map(A1 => l072_n_201, A2 => l072_n_149, ZN => l072_n_211);
  l072_g12457 : NR2D1BWP7T port map(A1 => l072_n_198, A2 => l072_n_113, ZN => l072_n_210);
  l072_g12458 : NR2D1BWP7T port map(A1 => l072_n_198, A2 => l072_n_114, ZN => l072_n_209);
  l072_g12459 : OAI21D0BWP7T port map(A1 => l072_n_131, A2 => l072_n_76, B => l072_n_199, ZN => l072_n_207);
  l072_g12460 : AOI21D0BWP7T port map(A1 => l072_n_143, A2 => l072_n_81, B => l072_n_204, ZN => l072_n_206);
  l072_g12461 : ND4D0BWP7T port map(A1 => l072_n_195, A2 => l072_n_190, A3 => l072_n_2, A4 => l072_n_182, ZN => l072_n_205);
  l072_g12462 : INVD0BWP7T port map(I => l072_n_203, ZN => l072_n_202);
  l072_g12463 : INVD0BWP7T port map(I => l072_n_201, ZN => l072_n_200);
  l072_g12464 : CKND2D1BWP7T port map(A1 => l072_n_193, A2 => l072_n_188, ZN => l072_n_204);
  l072_g12465 : NR2D1BWP7T port map(A1 => l072_n_194, A2 => l072_n_4, ZN => l072_n_203);
  l072_g12466 : NR2D1BWP7T port map(A1 => l072_n_194, A2 => l072_n_185, ZN => l072_n_201);
  l072_g12467 : OA31D1BWP7T port map(A1 => l072_n_120, A2 => l072_n_148, A3 => l072_n_175, B => l072_n_195, Z => l072_n_197);
  l072_g12468 : NR4D0BWP7T port map(A1 => l072_n_194, A2 => l072_n_173, A3 => l072_n_164, A4 => l072_n_43, ZN => l072_n_196);
  l072_g12469 : AOI21D0BWP7T port map(A1 => l072_n_2, A2 => l072_n_182, B => l072_n_194, ZN => l072_n_199);
  l072_g12470 : ND3D0BWP7T port map(A1 => l072_n_193, A2 => l072_n_176, A3 => l072_n_121, ZN => l072_n_198);
  l072_g12471 : INR2XD0BWP7T port map(A1 => l072_n_187, B1 => l072_n_192, ZN => l072_n_195);
  l072_g12472 : INVD1BWP7T port map(I => l072_n_194, ZN => l072_n_193);
  l072_g12473 : OAI221D0BWP7T port map(A1 => l072_n_174, A2 => l072_n_142, B1 => l072_n_29, B2 => l072_n_20, C => l072_n_191, ZN => l072_n_194);
  l072_g12474 : OAI221D0BWP7T port map(A1 => l072_n_185, A2 => l072_n_179, B1 => l072_n_171, B2 => l072_n_4, C => l072_n_181, ZN => l072_n_192);
  l072_g12475 : AOI221D0BWP7T port map(A1 => l072_n_8, A2 => x_enemy2(8), B1 => l072_n_51, B2 => l072_n_17, C => l072_n_186, ZN => l072_n_191);
  l072_g12476 : IAO21D0BWP7T port map(A1 => l072_n_4, A2 => l072_n_183, B => l072_n_189, ZN => l072_n_190);
  l072_g12477 : AOI21D0BWP7T port map(A1 => l072_n_183, A2 => l072_n_171, B => l072_n_185, ZN => l072_n_189);
  l072_g12478 : OAI22D0BWP7T port map(A1 => l072_n_4, A2 => l072_n_168, B1 => l072_n_185, B2 => l072_n_170, ZN => l072_n_188);
  l072_g12479 : IND2D1BWP7T port map(A1 => l072_n_4, B1 => l072_n_149, ZN => l072_n_187);
  l072_g12480 : AO21D0BWP7T port map(A1 => l072_n_20, A2 => l072_n_29, B => l072_n_180, Z => l072_n_186);
  l072_g12482 : NR3D0BWP7T port map(A1 => l072_n_163, A2 => l072_n_91, A3 => l072_n_64, ZN => l072_n_184);
  l072_g12483 : ND2D1BWP7T port map(A1 => l072_n_176, A2 => l072_n_119, ZN => l072_n_185);
  l072_g12485 : MOAI22D0BWP7T port map(A1 => l072_n_51, A2 => l072_n_17, B1 => l072_n_160, B2 => l072_n_142, ZN => l072_n_180);
  l072_g12486 : INR3D0BWP7T port map(A1 => l072_n_168, B1 => l072_n_166, B2 => l072_n_167, ZN => l072_n_183);
  l072_g12487 : ND4D0BWP7T port map(A1 => l072_n_0, A2 => l072_n_155, A3 => l072_n_146, A4 => l072_n_43, ZN => l072_n_182);
  l072_g12488 : IND3D1BWP7T port map(A1 => l072_n_148, B1 => l072_n_120, B2 => l072_n_177, ZN => l072_n_181);
  l072_g12489 : CKND1BWP7T port map(I => l072_n_178, ZN => l072_n_179);
  l072_g12490 : INVD0BWP7T port map(I => l072_n_176, ZN => l072_n_175);
  l072_g12491 : ND2D1BWP7T port map(A1 => l072_n_170, A2 => l072_n_165, ZN => l072_n_178);
  l072_g12492 : AOI211XD0BWP7T port map(A1 => l072_n_46, A2 => l072_n_30, B => l072_n_164, C => l072_n_101, ZN => l072_n_177);
  l072_g12493 : AOI211XD0BWP7T port map(A1 => l072_n_46, A2 => l072_n_24, B => l072_n_164, C => l072_n_100, ZN => l072_n_176);
  l072_g12494 : AOI221D0BWP7T port map(A1 => l072_n_107, A2 => l072_n_15, B1 => l072_n_49, B2 => l072_n_104, C => l072_n_159, ZN => l072_n_174);
  l072_g12495 : AOI22D0BWP7T port map(A1 => l072_n_0, A2 => y(4), B1 => l072_n_154, B2 => l072_n_41, ZN => l072_n_173);
  l072_g12496 : INR4D0BWP7T port map(A1 => l072_n_96, B1 => l072_n_94, B2 => l072_n_133, B3 => l072_n_147, ZN => l072_n_172);
  l072_g12497 : INVD0BWP7T port map(I => l072_n_170, ZN => l072_n_169);
  l072_g12498 : ND2D1BWP7T port map(A1 => l072_n_150, A2 => l072_n_113, ZN => l072_n_171);
  l072_g12499 : ND2D1BWP7T port map(A1 => l072_n_3, A2 => l072_n_113, ZN => l072_n_170);
  l072_g12500 : ND2D1BWP7T port map(A1 => l072_n_151, A2 => l072_n_114, ZN => l072_n_168);
  l072_g12501 : INR2D1BWP7T port map(A1 => l072_n_114, B1 => l072_n_158, ZN => l072_n_167);
  l072_g12502 : AN2D1BWP7T port map(A1 => l072_n_5, A2 => l072_n_113, Z => l072_n_166);
  l072_g12503 : ND2D1BWP7T port map(A1 => l072_n_152, A2 => l072_n_114, ZN => l072_n_165);
  l072_g12504 : IND4D0BWP7T port map(A1 => l072_n_71, B1 => l072_n_72, B2 => l072_n_102, B3 => l072_n_116, ZN => l072_n_163);
  l072_g12505 : ND4D0BWP7T port map(A1 => l072_n_129, A2 => l072_n_95, A3 => l072_n_70, A4 => l072_n_60, ZN => l072_n_162);
  l072_g12506 : IND4D0BWP7T port map(A1 => l072_n_76, B1 => l072_n_77, B2 => l072_n_70, B3 => l072_n_124, ZN => l072_n_161);
  l072_g12507 : OAI222D0BWP7T port map(A1 => l072_n_145, A2 => l072_n_138, B1 => l072_n_98, B2 => l072_n_137, C1 => l072_n_104, C2 => l072_n_105, ZN => l072_n_160);
  l072_g12508 : MOAI22D0BWP7T port map(A1 => l072_n_144, A2 => l072_n_136, B1 => l072_n_138, B2 => l072_n_106, ZN => l072_n_159);
  l072_g12509 : ND3D0BWP7T port map(A1 => l072_n_140, A2 => l072_n_146, A3 => l072_n_141, ZN => l072_n_164);
  l072_g12510 : OAI211D1BWP7T port map(A1 => l072_n_13, A2 => l072_n_56, B => l072_n_143, C => l072_n_89, ZN => l072_n_157);
  l072_g12511 : INR3D0BWP7T port map(A1 => l072_n_116, B1 => l072_n_93, B2 => l072_n_125, ZN => l072_n_156);
  l072_g12512 : AOI211D1BWP7T port map(A1 => l072_n_48, A2 => y(5), B => l072_n_123, C => l072_n_109, ZN => l072_n_155);
  l072_g12513 : NR3D0BWP7T port map(A1 => l072_n_134, A2 => l072_n_46, A3 => y(4), ZN => l072_n_154);
  l072_g12514 : AO211D0BWP7T port map(A1 => l072_n_59, A2 => l072_n_11, B => l072_n_147, C => l072_n_86, Z => l072_n_153);
  l072_g12515 : ND3D0BWP7T port map(A1 => l072_n_115, A2 => l072_n_110, A3 => l072_n_45, ZN => l072_n_158);
  l072_g12518 : NR3D0BWP7T port map(A1 => l072_n_117, A2 => l072_n_45, A3 => l072_n_47, ZN => l072_n_152);
  l072_g12520 : NR3D0BWP7T port map(A1 => l072_n_122, A2 => l072_n_115, A3 => l072_n_44, ZN => l072_n_151);
  l072_g12521 : AN4D1BWP7T port map(A1 => l072_n_115, A2 => l072_n_108, A3 => l072_n_1, A4 => l072_n_45, Z => l072_n_150);
  l072_g12522 : INR2D1BWP7T port map(A1 => l072_n_118, B1 => l072_n_135, ZN => l072_n_149);
  l072_g12523 : OR2D1BWP7T port map(A1 => l072_n_134, A2 => l072_n_41, Z => l072_n_148);
  l072_g12524 : ND2D1BWP7T port map(A1 => l072_n_132, A2 => l072_n_95, ZN => l072_n_147);
  l072_g12525 : AOI211XD0BWP7T port map(A1 => l072_n_53, A2 => l072_n_33, B => l072_n_90, C => l072_n_111, ZN => l072_n_146);
  l072_g12526 : CKND1BWP7T port map(I => l072_n_144, ZN => l072_n_145);
  l072_g12527 : AOI22D0BWP7T port map(A1 => l072_n_99, A2 => y(5), B1 => l072_n_83, B2 => y_enemy2(5), ZN => l072_n_141);
  l072_g12528 : NR2XD0BWP7T port map(A1 => l072_n_123, A2 => l072_n_109, ZN => l072_n_140);
  l072_g12529 : MAOI222D1BWP7T port map(A => l072_n_88, B => x(2), C => x_enemy2(2), ZN => l072_n_144);
  l072_g12530 : NR3D0BWP7T port map(A1 => l072_n_97, A2 => l072_n_91, A3 => l072_n_69, ZN => l072_n_143);
  l072_g12531 : OAI21D0BWP7T port map(A1 => l072_n_107, A2 => l072_n_14, B => l072_n_105, ZN => l072_n_142);
  l072_g12532 : CKND1BWP7T port map(I => l072_n_136, ZN => l072_n_137);
  l072_g12533 : INVD0BWP7T port map(I => l072_n_132, ZN => l072_n_131);
  l072_g12534 : AOI211XD0BWP7T port map(A1 => l072_n_59, A2 => l072_n_25, B => l072_n_97, C => l072_n_80, ZN => l072_n_130);
  l072_g12535 : OAI21D0BWP7T port map(A1 => l072_n_74, A2 => l072_n_58, B => draw_count6(1), ZN => l072_n_129);
  l072_g12536 : AOI221D0BWP7T port map(A1 => l072_n_58, A2 => l072_n_26, B1 => l072_n_62, B2 => draw_count6(0), C => l072_n_78, ZN => l072_n_128);
  l072_g12537 : AO221D0BWP7T port map(A1 => l072_n_66, A2 => l072_n_64, B1 => l072_n_67, B2 => l072_n_27, C => l072_n_94, Z => l072_n_127);
  l072_g12538 : OA211D0BWP7T port map(A1 => l072_n_25, A2 => l072_n_60, B => l072_n_102, C => l072_n_79, Z => l072_n_126);
  l072_g12539 : OAI211D1BWP7T port map(A1 => l072_n_11, A2 => l072_n_56, B => l072_n_81, C => l072_n_75, ZN => l072_n_125);
  l072_g12540 : AOI21D0BWP7T port map(A1 => l072_n_59, A2 => l072_n_26, B => l072_n_87, ZN => l072_n_124);
  l072_g12541 : AO21D0BWP7T port map(A1 => l072_n_67, A2 => l072_n_66, B => l072_n_94, Z => l072_n_139);
  l072_g12542 : OAI22D0BWP7T port map(A1 => l072_n_68, A2 => l072_n_16, B1 => l072_n_50, B2 => x(2), ZN => l072_n_138);
  l072_g12543 : IOA21D1BWP7T port map(A1 => l072_n_50, A2 => x(2), B => l072_n_106, ZN => l072_n_136);
  l072_g12544 : ND2D1BWP7T port map(A1 => l072_n_103, A2 => l072_n_42, ZN => l072_n_135);
  l072_g12545 : ND2D1BWP7T port map(A1 => l072_n_103, A2 => l072_n_84, ZN => l072_n_134);
  l072_g12546 : IND2D1BWP7T port map(A1 => l072_n_93, B1 => l072_n_70, ZN => l072_n_133);
  l072_g12547 : INR2XD0BWP7T port map(A1 => l072_n_60, B1 => l072_n_91, ZN => l072_n_132);
  l072_g12552 : OAI22D0BWP7T port map(A1 => l072_n_52, A2 => l072_n_28, B1 => l072_n_48, B2 => y(5), ZN => l072_n_123);
  l072_g12553 : MOAI22D0BWP7T port map(A1 => l072_n_60, A2 => draw_count6(1), B1 => l072_n_74, B2 => l072_n_66, ZN => l072_n_112);
  l072_g12554 : MOAI22D0BWP7T port map(A1 => l072_n_19, A2 => y(9), B1 => l072_n_19, B2 => y(9), ZN => l072_n_111);
  l072_g12555 : MAOI22D0BWP7T port map(A1 => l072_n_84, A2 => l072_n_34, B1 => l072_n_84, B2 => l072_n_34, ZN => l072_n_122);
  l072_g12556 : MAOI22D0BWP7T port map(A1 => l072_n_43, A2 => l072_n_35, B1 => l072_n_43, B2 => l072_n_35, ZN => l072_n_121);
  l072_g12557 : MAOI22D0BWP7T port map(A1 => l072_n_43, A2 => y(3), B1 => l072_n_43, B2 => y(3), ZN => l072_n_120);
  l072_g12558 : MOAI22D0BWP7T port map(A1 => l072_n_43, A2 => l072_n_18, B1 => l072_n_43, B2 => l072_n_18, ZN => l072_n_119);
  l072_g12559 : MAOI22D0BWP7T port map(A1 => l072_n_82, A2 => y(2), B1 => l072_n_82, B2 => y(2), ZN => l072_n_118);
  l072_g12560 : ND2D1BWP7T port map(A1 => l072_n_108, A2 => l072_n_1, ZN => l072_n_110);
  l072_g12561 : MAOI22D0BWP7T port map(A1 => l072_n_42, A2 => y(1), B1 => l072_n_42, B2 => y(1), ZN => l072_n_117);
  l072_g12562 : INR3D0BWP7T port map(A1 => l072_n_79, B1 => l072_n_62, B2 => l072_n_78, ZN => l072_n_116);
  l072_g12563 : MOAI22D0BWP7T port map(A1 => l072_n_47, A2 => y(0), B1 => l072_n_47, B2 => y(0), ZN => l072_n_115);
  l072_g12564 : MAOI22D0BWP7T port map(A1 => l072_n_41, A2 => l072_n_21, B1 => l072_n_41, B2 => l072_n_21, ZN => l072_n_114);
  l072_g12565 : MOAI22D0BWP7T port map(A1 => l072_n_41, A2 => l072_n_23, B1 => l072_n_41, B2 => l072_n_23, ZN => l072_n_113);
  l072_g12566 : NR2XD0BWP7T port map(A1 => l072_n_46, A2 => l072_n_30, ZN => l072_n_101);
  l072_g12567 : NR2XD0BWP7T port map(A1 => l072_n_46, A2 => l072_n_24, ZN => l072_n_100);
  l072_g12569 : CKAN2D1BWP7T port map(A1 => l072_n_52, A2 => l072_n_28, Z => l072_n_109);
  l072_g12570 : ND2D1BWP7T port map(A1 => l072_n_42, A2 => l072_n_31, ZN => l072_n_108);
  l072_g12571 : NR2D1BWP7T port map(A1 => l072_n_83, A2 => y_enemy2(5), ZN => l072_n_99);
  l072_g12572 : CKAN2D1BWP7T port map(A1 => l072_n_49, A2 => l072_n_38, Z => l072_n_107);
  l072_g12573 : ND2D1BWP7T port map(A1 => l072_n_68, A2 => l072_n_16, ZN => l072_n_106);
  l072_g12574 : OR2D1BWP7T port map(A1 => l072_n_49, A2 => l072_n_15, Z => l072_n_105);
  l072_g12575 : NR2XD0BWP7T port map(A1 => l072_n_68, A2 => l072_n_16, ZN => l072_n_98);
  l072_g12576 : CKAN2D1BWP7T port map(A1 => l072_n_14, A2 => l072_n_38, Z => l072_n_104);
  l072_g12577 : INR2D1BWP7T port map(A1 => l072_n_47, B1 => l072_n_45, ZN => l072_n_103);
  l072_g12578 : NR2XD0BWP7T port map(A1 => l072_n_73, A2 => l072_n_80, ZN => l072_n_102);
  l072_g12579 : NR2D0BWP7T port map(A1 => l072_n_53, A2 => l072_n_33, ZN => l072_n_90);
  l072_g12580 : AOI22D0BWP7T port map(A1 => l072_n_59, A2 => l072_n_12, B1 => l072_n_62, B2 => l072_n_25, ZN => l072_n_89);
  l072_g12581 : AOI22D0BWP7T port map(A1 => l072_n_54, A2 => x(0), B1 => x(1), B2 => l072_n_9, ZN => l072_n_88);
  l072_g12582 : AOI21D0BWP7T port map(A1 => l072_n_57, A2 => l072_n_60, B => draw_count6(1), ZN => l072_n_87);
  l072_g12583 : OA21D0BWP7T port map(A1 => l072_n_58, A2 => l072_n_55, B => l072_n_25, Z => l072_n_86);
  l072_g12584 : AOI21D0BWP7T port map(A1 => l072_n_58, A2 => l072_n_25, B => l072_n_63, ZN => l072_n_85);
  l072_g12585 : OAI21D0BWP7T port map(A1 => l072_n_56, A2 => draw_count6(1), B => l072_n_75, ZN => l072_n_97);
  l072_g12586 : AOI21D0BWP7T port map(A1 => l072_n_62, A2 => l072_n_11, B => l072_n_59, ZN => l072_n_96);
  l072_g12587 : OAI21D0BWP7T port map(A1 => l072_n_63, A2 => l072_n_55, B => l072_n_12, ZN => l072_n_95);
  l072_g12588 : MOAI22D0BWP7T port map(A1 => l072_n_65, A2 => l072_n_26, B1 => l072_n_67, B2 => l072_n_12, ZN => l072_n_94);
  l072_g12589 : AO21D0BWP7T port map(A1 => l072_n_64, A2 => l072_n_26, B => l072_n_73, Z => l072_n_93);
  l072_g12590 : IOA21D1BWP7T port map(A1 => l072_n_58, A2 => l072_n_11, B => l072_n_77, ZN => l072_n_92);
  l072_g12591 : OAI22D0BWP7T port map(A1 => l072_n_57, A2 => l072_n_11, B1 => l072_n_60, B2 => l072_n_26, ZN => l072_n_91);
  l072_g12592 : INVD1BWP7T port map(I => l072_n_42, ZN => l072_n_84);
  l072_g12594 : INVD0BWP7T port map(I => l072_n_48, ZN => l072_n_83);
  l072_g12595 : INVD0BWP7T port map(I => l072_n_41, ZN => l072_n_82);
  l072_g12596 : ND2D1BWP7T port map(A1 => l072_n_59, A2 => draw_count6(1), ZN => l072_n_81);
  l072_g12597 : NR2D1BWP7T port map(A1 => l072_n_65, A2 => draw_count6(1), ZN => l072_n_80);
  l072_g12598 : IND2D0BWP7T port map(A1 => l072_n_13, B1 => l072_n_63, ZN => l072_n_79);
  l072_g12599 : INR2D1BWP7T port map(A1 => l072_n_59, B1 => draw_count6(1), ZN => l072_n_78);
  l072_g12600 : CKND2D0BWP7T port map(A1 => l072_n_63, A2 => l072_n_12, ZN => l072_n_77);
  l072_g12601 : NR2D0BWP7T port map(A1 => l072_n_56, A2 => l072_n_6, ZN => l072_n_76);
  l072_g12602 : NR2D0BWP7T port map(A1 => l072_n_60, A2 => l072_n_13, ZN => l072_n_69);
  l072_g12603 : CKND2D1BWP7T port map(A1 => l072_n_58, A2 => l072_n_66, ZN => l072_n_75);
  l072_g12604 : IND2D1BWP7T port map(A1 => l072_n_59, B1 => l072_n_61, ZN => l072_n_74);
  l072_g12605 : AN2D0BWP7T port map(A1 => l072_n_63, A2 => l072_n_25, Z => l072_n_73);
  l072_g12606 : ND2D1BWP7T port map(A1 => l072_n_55, A2 => l072_n_11, ZN => l072_n_72);
  l072_g12607 : INR2D1BWP7T port map(A1 => l072_n_27, B1 => l072_n_57, ZN => l072_n_71);
  l072_g12608 : ND2D1BWP7T port map(A1 => l072_n_63, A2 => l072_n_66, ZN => l072_n_70);
  l072_g12609 : INVD1BWP7T port map(I => l072_n_65, ZN => l072_n_64);
  l072_g12610 : INVD1BWP7T port map(I => l072_n_62, ZN => l072_n_61);
  l072_g12611 : INVD0BWP7T port map(I => l072_n_58, ZN => l072_n_57);
  l072_g12612 : INVD1BWP7T port map(I => l072_n_56, ZN => l072_n_55);
  l072_g12613 : IAO21D0BWP7T port map(A1 => x(1), A2 => l072_n_9, B => x_enemy2(0), ZN => l072_n_54);
  l072_g12614 : AO21D0BWP7T port map(A1 => x(4), A2 => l072_n_10, B => l072_n_14, Z => l072_n_68);
  l072_g12615 : INR2D1BWP7T port map(A1 => draw_count6(3), B1 => l072_n_32, ZN => l072_n_67);
  l072_g12616 : IND2D1BWP7T port map(A1 => l072_n_27, B1 => l072_n_13, ZN => l072_n_66);
  l072_g12617 : ND2D1BWP7T port map(A1 => l072_n_39, A2 => draw_count6(3), ZN => l072_n_65);
  l072_g12618 : NR2D1BWP7T port map(A1 => l072_n_32, A2 => draw_count6(3), ZN => l072_n_63);
  l072_g12619 : INR2D1BWP7T port map(A1 => l072_n_22, B1 => draw_count6(3), ZN => l072_n_62);
  l072_g12620 : ND2D1BWP7T port map(A1 => l072_n_36, A2 => draw_count6(3), ZN => l072_n_60);
  l072_g12621 : NR2D1BWP7T port map(A1 => l072_n_37, A2 => draw_count6(3), ZN => l072_n_59);
  l072_g12622 : NR2D1BWP7T port map(A1 => l072_n_40, A2 => draw_count6(3), ZN => l072_n_58);
  l072_g12623 : ND2D1BWP7T port map(A1 => l072_n_22, A2 => draw_count6(3), ZN => l072_n_56);
  l072_g12625 : INVD0BWP7T port map(I => l072_n_45, ZN => l072_n_44);
  l072_g12626 : MOAI22D0BWP7T port map(A1 => y(8), A2 => y_enemy2(8), B1 => y(8), B2 => y_enemy2(8), ZN => l072_n_53);
  l072_g12627 : MAOI22D0BWP7T port map(A1 => y(7), A2 => y_enemy2(7), B1 => y(7), B2 => y_enemy2(7), ZN => l072_n_52);
  l072_g12628 : MOAI22D0BWP7T port map(A1 => x(7), A2 => x_enemy2(7), B1 => x(7), B2 => x_enemy2(7), ZN => l072_n_51);
  l072_g12629 : MAOI22D0BWP7T port map(A1 => x(3), A2 => x_enemy2(3), B1 => x(3), B2 => x_enemy2(3), ZN => l072_n_50);
  l072_g12630 : MAOI22D0BWP7T port map(A1 => x(6), A2 => x_enemy2(6), B1 => x(6), B2 => x_enemy2(6), ZN => l072_n_49);
  l072_g12631 : OAI21D0BWP7T port map(A1 => l072_n_7, A2 => y_enemy2(6), B => l072_n_28, ZN => l072_n_48);
  l072_g12632 : MOAI22D0BWP7T port map(A1 => y(1), A2 => y_enemy2(1), B1 => y(1), B2 => y_enemy2(1), ZN => l072_n_47);
  l072_g12633 : MAOI22D0BWP7T port map(A1 => y(5), A2 => y_enemy2(5), B1 => y(5), B2 => y_enemy2(5), ZN => l072_n_46);
  l072_g12634 : MAOI22D0BWP7T port map(A1 => y(0), A2 => y_enemy2(0), B1 => y(0), B2 => y_enemy2(0), ZN => l072_n_45);
  l072_g12635 : MOAI22D0BWP7T port map(A1 => y(4), A2 => y_enemy2(4), B1 => y(4), B2 => y_enemy2(4), ZN => l072_n_43);
  l072_g12636 : MAOI22D0BWP7T port map(A1 => y(2), A2 => y_enemy2(2), B1 => y(2), B2 => y_enemy2(2), ZN => l072_n_42);
  l072_g12637 : MOAI22D0BWP7T port map(A1 => y(3), A2 => y_enemy2(3), B1 => y(3), B2 => y_enemy2(3), ZN => l072_n_41);
  l072_g12638 : CKND1BWP7T port map(I => l072_n_39, ZN => l072_n_40);
  l072_g12639 : CKND1BWP7T port map(I => l072_n_36, ZN => l072_n_37);
  l072_g12640 : INVD1BWP7T port map(I => l072_n_26, ZN => l072_n_25);
  l072_g12641 : INR2D1BWP7T port map(A1 => draw_count6(4), B1 => draw_count6(2), ZN => l072_n_39);
  l072_g12642 : IND2D1BWP7T port map(A1 => x_enemy2(5), B1 => x(5), ZN => l072_n_38);
  l072_g12643 : INR2D1BWP7T port map(A1 => draw_count6(2), B1 => draw_count6(4), ZN => l072_n_36);
  l072_g12644 : IND2D0BWP7T port map(A1 => y_enemy2(3), B1 => y(3), ZN => l072_n_35);
  l072_g12645 : IND2D1BWP7T port map(A1 => y_enemy2(1), B1 => y(1), ZN => l072_n_34);
  l072_g12646 : INR2XD0BWP7T port map(A1 => y_enemy2(7), B1 => y(7), ZN => l072_n_33);
  l072_g12647 : ND2D1BWP7T port map(A1 => draw_count6(2), A2 => draw_count6(4), ZN => l072_n_32);
  l072_g12648 : IND2D1BWP7T port map(A1 => y(1), B1 => y_enemy2(1), ZN => l072_n_31);
  l072_g12649 : IND2D0BWP7T port map(A1 => y_enemy2(4), B1 => y(4), ZN => l072_n_30);
  l072_g12650 : IND2D1BWP7T port map(A1 => x(7), B1 => x_enemy2(7), ZN => l072_n_29);
  l072_g12651 : ND2D1BWP7T port map(A1 => l072_n_7, A2 => y_enemy2(6), ZN => l072_n_28);
  l072_g12652 : INR2D1BWP7T port map(A1 => draw_count6(0), B1 => draw_count6(1), ZN => l072_n_27);
  l072_g12653 : CKND2D1BWP7T port map(A1 => draw_count6(1), A2 => draw_count6(0), ZN => l072_n_26);
  l072_g12654 : INVD1BWP7T port map(I => l072_n_12, ZN => l072_n_11);
  l072_g12655 : INR2XD0BWP7T port map(A1 => y_enemy2(4), B1 => y(4), ZN => l072_n_24);
  l072_g12656 : IND2D1BWP7T port map(A1 => y(2), B1 => y_enemy2(2), ZN => l072_n_23);
  l072_g12657 : NR2D0BWP7T port map(A1 => draw_count6(2), A2 => draw_count6(4), ZN => l072_n_22);
  l072_g12658 : IND2D1BWP7T port map(A1 => y_enemy2(2), B1 => y(2), ZN => l072_n_21);
  l072_g12659 : NR2D1BWP7T port map(A1 => l072_n_8, A2 => x_enemy2(8), ZN => l072_n_20);
  l072_g12660 : IND2D1BWP7T port map(A1 => y(8), B1 => y_enemy2(8), ZN => l072_n_19);
  l072_g12661 : IND2D1BWP7T port map(A1 => y(3), B1 => y_enemy2(3), ZN => l072_n_18);
  l072_g12662 : IND2D1BWP7T port map(A1 => x_enemy2(6), B1 => x(6), ZN => l072_n_17);
  l072_g12663 : IND2D1BWP7T port map(A1 => x(3), B1 => x_enemy2(3), ZN => l072_n_16);
  l072_g12664 : INR2XD0BWP7T port map(A1 => x_enemy2(5), B1 => x(5), ZN => l072_n_15);
  l072_g12665 : NR2D1BWP7T port map(A1 => x(4), A2 => l072_n_10, ZN => l072_n_14);
  l072_g12666 : IND2D1BWP7T port map(A1 => draw_count6(0), B1 => draw_count6(1), ZN => l072_n_13);
  l072_g12667 : NR2D0BWP7T port map(A1 => draw_count6(1), A2 => draw_count6(0), ZN => l072_n_12);
  l072_g12668 : INVD0BWP7T port map(I => x_enemy2(4), ZN => l072_n_10);
  l072_g12669 : INVD0BWP7T port map(I => x_enemy2(1), ZN => l072_n_9);
  l072_g12670 : CKND1BWP7T port map(I => x(8), ZN => l072_n_8);
  l072_g12671 : INVD1BWP7T port map(I => y(6), ZN => l072_n_7);
  l072_g12672 : INVD0BWP7T port map(I => draw_count6(1), ZN => l072_n_6);
  l072_g2 : INR3D0BWP7T port map(A1 => l072_n_122, B1 => l072_n_115, B2 => l072_n_44, ZN => l072_n_5);
  l072_g12673 : IND2D1BWP7T port map(A1 => l072_n_119, B1 => l072_n_177, ZN => l072_n_4);
  l072_g12674 : INR3D0BWP7T port map(A1 => l072_n_117, B1 => l072_n_45, B2 => l072_n_47, ZN => l072_n_3);
  l072_g12675 : IIND4D0BWP7T port map(A1 => l072_n_121, A2 => l072_n_113, B1 => l072_n_150, B2 => l072_n_177, ZN => l072_n_2);
  l072_g12676 : IND2D1BWP7T port map(A1 => l072_n_31, B1 => l072_n_84, ZN => l072_n_1);
  l072_g12677 : INR3D0BWP7T port map(A1 => l072_n_46, B1 => l072_n_134, B2 => l072_n_82, ZN => l072_n_0);
  l01_count_reg_8 : DFQD1BWP7T port map(CP => clk, D => l01_n_31, Q => x(8));
  l01_g608 : AO211D0BWP7T port map(A1 => l01_n_23, A2 => x(8), B => l01_n_28, C => reset, Z => l01_n_31);
  l01_g609 : AO211D0BWP7T port map(A1 => l01_n_18, A2 => x(7), B => l01_n_27, C => reset, Z => l01_n_30);
  l01_g611 : AO211D0BWP7T port map(A1 => l01_n_21, A2 => x(6), B => l01_n_26, C => reset, Z => l01_n_29);
  l01_g612 : NR4D0BWP7T port map(A1 => l01_n_21, A2 => l01_n_0, A3 => l01_n_1, A4 => x(8), ZN => l01_n_28);
  l01_g613 : OAI32D0BWP7T port map(A1 => x(7), A2 => l01_n_1, A3 => l01_n_21, B1 => l01_n_7, B2 => l01_n_5, ZN => l01_n_27);
  l01_count_reg_5 : DFQD1BWP7T port map(CP => clk, D => l01_n_25, Q => x(5));
  l01_g616 : NR2D0BWP7T port map(A1 => l01_n_21, A2 => x(6), ZN => l01_n_26);
  l01_g617 : AO211D0BWP7T port map(A1 => l01_n_19, A2 => x(5), B => l01_n_22, C => reset, Z => l01_n_25);
  l01_g618 : AO211D0BWP7T port map(A1 => l01_n_16, A2 => x(4), B => l01_n_20, C => reset, Z => l01_n_24);
  l01_g619 : AO211D0BWP7T port map(A1 => l01_n_1, A2 => x(5), B => l01_n_18, C => l01_n_0, Z => l01_n_23);
  l01_g620 : NR2D0BWP7T port map(A1 => l01_n_19, A2 => x(5), ZN => l01_n_22);
  l01_count_reg_3 : DFQD1BWP7T port map(CP => clk, D => l01_n_17, Q => x(3));
  l01_g622 : AOI211D1BWP7T port map(A1 => l01_n_6, A2 => l01_n_7, B => l01_n_16, C => x(4), ZN => l01_n_20);
  l01_g623 : IND2D1BWP7T port map(A1 => l01_n_19, B1 => x(5), ZN => l01_n_21);
  l01_g624 : IND2D1BWP7T port map(A1 => l01_n_16, B1 => x(4), ZN => l01_n_19);
  l01_g625 : AO211D0BWP7T port map(A1 => l01_n_13, A2 => x(3), B => l01_n_15, C => reset, Z => l01_n_17);
  l01_g626 : OR2D1BWP7T port map(A1 => l01_n_10, A2 => l01_n_16, Z => l01_n_18);
  l01_count_reg_2 : DFQD1BWP7T port map(CP => clk, D => l01_n_14, Q => x(2));
  l01_g628 : IND2D1BWP7T port map(A1 => l01_n_13, B1 => x(3), ZN => l01_n_16);
  l01_g629 : NR2D0BWP7T port map(A1 => l01_n_13, A2 => x(3), ZN => l01_n_15);
  l01_g630 : AO211D0BWP7T port map(A1 => l01_n_9, A2 => x(2), B => l01_n_12, C => reset, Z => l01_n_14);
  l01_count_reg_1 : DFQD1BWP7T port map(CP => clk, D => l01_n_11, Q => x(1));
  l01_g632 : IND2D1BWP7T port map(A1 => l01_n_9, B1 => x(2), ZN => l01_n_13);
  l01_g633 : NR2D0BWP7T port map(A1 => l01_n_9, A2 => x(2), ZN => l01_n_12);
  l01_g634 : AO211D0BWP7T port map(A1 => l01_n_3, A2 => x(1), B => l01_n_8, C => reset, Z => l01_n_11);
  l01_g635 : OAI222D0BWP7T port map(A1 => l01_n_2, A2 => x(6), B1 => x(5), B2 => l01_n_1, C1 => x(4), C2 => l01_n_1, ZN => l01_n_10);
  l01_g637 : NR2D0BWP7T port map(A1 => l01_n_3, A2 => x(1), ZN => l01_n_8);
  l01_g638 : ND2D1BWP7T port map(A1 => x(1), A2 => x(0), ZN => l01_n_9);
  l01_g639 : CKND1BWP7T port map(I => l01_n_5, ZN => l01_n_6);
  l01_g640 : IND2D1BWP7T port map(A1 => reset, B1 => x(0), ZN => l01_n_4);
  l01_g641 : INR2XD0BWP7T port map(A1 => x(8), B1 => x(5), ZN => l01_n_7);
  l01_g642 : ND2D1BWP7T port map(A1 => l01_n_1, A2 => x(7), ZN => l01_n_5);
  l01_count_reg_7 : DFD1BWP7T port map(CP => clk, D => l01_n_30, Q => x(7), QN => l01_n_0);
  l01_count_reg_0 : DFD1BWP7T port map(CP => clk, D => l01_n_4, Q => x(0), QN => l01_n_3);
  l01_count_reg_4 : DFD1BWP7T port map(CP => clk, D => l01_n_24, Q => x(4), QN => l01_n_2);
  l01_count_reg_6 : DFD1BWP7T port map(CP => clk, D => l01_n_29, Q => x(6), QN => l01_n_1);
  l073_g12395 : OAI221D0BWP7T port map(A1 => l073_n_222, A2 => l073_n_184, B1 => l073_n_156, B2 => l073_n_225, C => l073_n_246, ZN => r7);
  l073_g12396 : NR4D0BWP7T port map(A1 => l073_n_245, A2 => l073_n_235, A3 => l073_n_229, A4 => l073_n_206, ZN => l073_n_246);
  l073_g12397 : IND4D0BWP7T port map(A1 => l073_n_233, B1 => l073_n_228, B2 => l073_n_234, B3 => l073_n_242, ZN => l073_n_245);
  l073_g12398 : AO211D0BWP7T port map(A1 => l073_n_218, A2 => l073_n_92, B => l073_n_243, C => l073_n_241, Z => g7);
  l073_g12399 : OAI211D1BWP7T port map(A1 => l073_n_126, A2 => l073_n_222, B => l073_n_239, C => l073_n_231, ZN => l073_n_243);
  l073_g12400 : MAOI22D0BWP7T port map(A1 => l073_n_215, A2 => l073_n_162, B1 => l073_n_236, B2 => l073_n_194, ZN => l073_n_242);
  l073_g12401 : AO221D0BWP7T port map(A1 => l073_n_215, A2 => l073_n_139, B1 => l073_n_212, B2 => l073_n_127, C => l073_n_237, Z => l073_n_241);
  l073_g12402 : OAI32D1BWP7T port map(A1 => l073_n_25, A2 => l073_n_61, A3 => l073_n_222, B1 => l073_n_96, B2 => l073_n_224, ZN => b7);
  l073_g12403 : AOI211XD0BWP7T port map(A1 => l073_n_199, A2 => l073_n_71, B => l073_n_232, C => l073_n_226, ZN => l073_n_239);
  l073_g12404 : ND3D0BWP7T port map(A1 => l073_n_220, A2 => l073_n_211, A3 => l073_n_198, ZN => enable7);
  l073_g12405 : OAI211D1BWP7T port map(A1 => l073_n_85, A2 => l073_n_204, B => l073_n_219, C => l073_n_227, ZN => l073_n_237);
  l073_g12406 : ND4D0BWP7T port map(A1 => l073_n_216, A2 => l073_n_187, A3 => l073_n_181, A4 => l073_n_165, ZN => l073_n_236);
  l073_g12407 : OAI211D1BWP7T port map(A1 => l073_n_172, A2 => l073_n_224, B => l073_n_221, C => l073_n_207, ZN => l073_n_235);
  l073_g12408 : AOI22D0BWP7T port map(A1 => l073_n_212, A2 => l073_n_157, B1 => l073_n_217, B2 => l073_n_161, ZN => l073_n_234);
  l073_g12409 : AOI31D0BWP7T port map(A1 => l073_n_130, A2 => l073_n_132, A3 => l073_n_61, B => l073_n_230, ZN => l073_n_233);
  l073_g12410 : AOI21D0BWP7T port map(A1 => l073_n_132, A2 => l073_n_72, B => l073_n_225, ZN => l073_n_232);
  l073_g12411 : OAI21D0BWP7T port map(A1 => l073_n_133, A2 => l073_n_92, B => l073_n_223, ZN => l073_n_231);
  l073_g12412 : AOI21D0BWP7T port map(A1 => l073_n_210, A2 => l073_n_150, B => l073_n_196, ZN => l073_n_230);
  l073_g12413 : IAO21D0BWP7T port map(A1 => l073_n_153, A2 => l073_n_71, B => l073_n_213, ZN => l073_n_229);
  l073_g12414 : OAI31D0BWP7T port map(A1 => l073_n_76, A2 => l073_n_92, A3 => l073_n_112, B => l073_n_214, ZN => l073_n_228);
  l073_g12415 : OAI21D0BWP7T port map(A1 => l073_n_133, A2 => l073_n_139, B => l073_n_214, ZN => l073_n_227);
  l073_g12416 : AOI21D0BWP7T port map(A1 => l073_n_102, A2 => l073_n_70, B => l073_n_213, ZN => l073_n_226);
  l073_g12417 : INVD0BWP7T port map(I => l073_n_223, ZN => l073_n_224);
  l073_g12418 : OAI21D0BWP7T port map(A1 => l073_n_91, A2 => l073_n_55, B => l073_n_218, ZN => l073_n_221);
  l073_g12419 : AOI22D0BWP7T port map(A1 => l073_n_205, A2 => l073_n_193, B1 => l073_n_203, B2 => l073_n_178, ZN => l073_n_220);
  l073_g12420 : OAI21D0BWP7T port map(A1 => l073_n_93, A2 => l073_n_64, B => l073_n_217, ZN => l073_n_219);
  l073_g12421 : AOI22D0BWP7T port map(A1 => l073_n_209, A2 => l073_n_151, B1 => l073_n_210, B2 => l073_n_3, ZN => l073_n_225);
  l073_g12422 : OAI32D1BWP7T port map(A1 => l073_n_118, A2 => l073_n_135, A3 => l073_n_198, B1 => l073_n_158, B2 => l073_n_208, ZN => l073_n_223);
  l073_g12423 : AOI22D0BWP7T port map(A1 => l073_n_210, A2 => l073_n_5, B1 => l073_n_209, B2 => l073_n_152, ZN => l073_n_222);
  l073_g12424 : AOI211D1BWP7T port map(A1 => l073_n_128, A2 => l073_n_56, B => l073_n_197, C => l073_n_188, ZN => l073_n_216);
  l073_g12425 : OAI22D0BWP7T port map(A1 => l073_n_200, A2 => l073_n_171, B1 => l073_n_194, B2 => l073_n_181, ZN => l073_n_218);
  l073_g12426 : IOA21D1BWP7T port map(A1 => l073_n_203, A2 => l073_n_167, B => l073_n_211, ZN => l073_n_217);
  l073_g12427 : MOAI22D0BWP7T port map(A1 => l073_n_200, A2 => l073_n_165, B1 => l073_n_203, B2 => l073_n_166, ZN => l073_n_215);
  l073_g12428 : MOAI22D0BWP7T port map(A1 => l073_n_200, A2 => l073_n_168, B1 => l073_n_203, B2 => l073_n_169, ZN => l073_n_214);
  l073_g12429 : MAOI22D0BWP7T port map(A1 => l073_n_201, A2 => l073_n_166, B1 => l073_n_202, B2 => l073_n_165, ZN => l073_n_213);
  l073_g12430 : MOAI22D0BWP7T port map(A1 => l073_n_194, A2 => l073_n_187, B1 => l073_n_201, B2 => l073_n_167, ZN => l073_n_212);
  l073_g12431 : INVD0BWP7T port map(I => l073_n_209, ZN => l073_n_208);
  l073_g12432 : ND2D1BWP7T port map(A1 => l073_n_201, A2 => l073_n_149, ZN => l073_n_211);
  l073_g12433 : NR2D1BWP7T port map(A1 => l073_n_198, A2 => l073_n_113, ZN => l073_n_210);
  l073_g12434 : NR2D1BWP7T port map(A1 => l073_n_198, A2 => l073_n_114, ZN => l073_n_209);
  l073_g12435 : OAI21D0BWP7T port map(A1 => l073_n_131, A2 => l073_n_76, B => l073_n_199, ZN => l073_n_207);
  l073_g12436 : AOI21D0BWP7T port map(A1 => l073_n_143, A2 => l073_n_81, B => l073_n_204, ZN => l073_n_206);
  l073_g12437 : ND4D0BWP7T port map(A1 => l073_n_195, A2 => l073_n_190, A3 => l073_n_2, A4 => l073_n_182, ZN => l073_n_205);
  l073_g12438 : INVD0BWP7T port map(I => l073_n_203, ZN => l073_n_202);
  l073_g12439 : INVD0BWP7T port map(I => l073_n_201, ZN => l073_n_200);
  l073_g12440 : CKND2D1BWP7T port map(A1 => l073_n_193, A2 => l073_n_188, ZN => l073_n_204);
  l073_g12441 : NR2D1BWP7T port map(A1 => l073_n_194, A2 => l073_n_4, ZN => l073_n_203);
  l073_g12442 : NR2D1BWP7T port map(A1 => l073_n_194, A2 => l073_n_185, ZN => l073_n_201);
  l073_g12443 : OA31D1BWP7T port map(A1 => l073_n_120, A2 => l073_n_148, A3 => l073_n_175, B => l073_n_195, Z => l073_n_197);
  l073_g12444 : NR4D0BWP7T port map(A1 => l073_n_194, A2 => l073_n_173, A3 => l073_n_164, A4 => l073_n_43, ZN => l073_n_196);
  l073_g12445 : AOI21D0BWP7T port map(A1 => l073_n_2, A2 => l073_n_182, B => l073_n_194, ZN => l073_n_199);
  l073_g12446 : ND3D0BWP7T port map(A1 => l073_n_193, A2 => l073_n_176, A3 => l073_n_121, ZN => l073_n_198);
  l073_g12447 : INR2XD0BWP7T port map(A1 => l073_n_187, B1 => l073_n_192, ZN => l073_n_195);
  l073_g12448 : INVD1BWP7T port map(I => l073_n_194, ZN => l073_n_193);
  l073_g12449 : OAI221D0BWP7T port map(A1 => l073_n_174, A2 => l073_n_142, B1 => l073_n_29, B2 => l073_n_20, C => l073_n_191, ZN => l073_n_194);
  l073_g12450 : OAI221D0BWP7T port map(A1 => l073_n_185, A2 => l073_n_179, B1 => l073_n_171, B2 => l073_n_4, C => l073_n_181, ZN => l073_n_192);
  l073_g12451 : AOI221D0BWP7T port map(A1 => l073_n_8, A2 => x_enemy3(8), B1 => l073_n_51, B2 => l073_n_17, C => l073_n_186, ZN => l073_n_191);
  l073_g12452 : IAO21D0BWP7T port map(A1 => l073_n_4, A2 => l073_n_183, B => l073_n_189, ZN => l073_n_190);
  l073_g12453 : AOI21D0BWP7T port map(A1 => l073_n_183, A2 => l073_n_171, B => l073_n_185, ZN => l073_n_189);
  l073_g12454 : OAI22D0BWP7T port map(A1 => l073_n_4, A2 => l073_n_168, B1 => l073_n_185, B2 => l073_n_170, ZN => l073_n_188);
  l073_g12455 : IND2D1BWP7T port map(A1 => l073_n_4, B1 => l073_n_149, ZN => l073_n_187);
  l073_g12456 : AO21D0BWP7T port map(A1 => l073_n_20, A2 => l073_n_29, B => l073_n_180, Z => l073_n_186);
  l073_g12458 : NR3D0BWP7T port map(A1 => l073_n_163, A2 => l073_n_91, A3 => l073_n_64, ZN => l073_n_184);
  l073_g12459 : ND2D1BWP7T port map(A1 => l073_n_176, A2 => l073_n_119, ZN => l073_n_185);
  l073_g12461 : MOAI22D0BWP7T port map(A1 => l073_n_51, A2 => l073_n_17, B1 => l073_n_160, B2 => l073_n_142, ZN => l073_n_180);
  l073_g12462 : INR3D0BWP7T port map(A1 => l073_n_168, B1 => l073_n_166, B2 => l073_n_167, ZN => l073_n_183);
  l073_g12463 : ND4D0BWP7T port map(A1 => l073_n_0, A2 => l073_n_155, A3 => l073_n_146, A4 => l073_n_43, ZN => l073_n_182);
  l073_g12464 : IND3D1BWP7T port map(A1 => l073_n_148, B1 => l073_n_120, B2 => l073_n_177, ZN => l073_n_181);
  l073_g12465 : CKND1BWP7T port map(I => l073_n_178, ZN => l073_n_179);
  l073_g12466 : INVD0BWP7T port map(I => l073_n_176, ZN => l073_n_175);
  l073_g12467 : ND2D1BWP7T port map(A1 => l073_n_170, A2 => l073_n_165, ZN => l073_n_178);
  l073_g12468 : AOI211XD0BWP7T port map(A1 => l073_n_46, A2 => l073_n_30, B => l073_n_164, C => l073_n_101, ZN => l073_n_177);
  l073_g12469 : AOI211XD0BWP7T port map(A1 => l073_n_46, A2 => l073_n_24, B => l073_n_164, C => l073_n_100, ZN => l073_n_176);
  l073_g12470 : AOI221D0BWP7T port map(A1 => l073_n_107, A2 => l073_n_15, B1 => l073_n_49, B2 => l073_n_104, C => l073_n_159, ZN => l073_n_174);
  l073_g12471 : AOI22D0BWP7T port map(A1 => l073_n_0, A2 => y(4), B1 => l073_n_154, B2 => l073_n_41, ZN => l073_n_173);
  l073_g12472 : INR4D0BWP7T port map(A1 => l073_n_96, B1 => l073_n_94, B2 => l073_n_133, B3 => l073_n_147, ZN => l073_n_172);
  l073_g12473 : INVD0BWP7T port map(I => l073_n_170, ZN => l073_n_169);
  l073_g12474 : ND2D1BWP7T port map(A1 => l073_n_150, A2 => l073_n_113, ZN => l073_n_171);
  l073_g12475 : ND2D1BWP7T port map(A1 => l073_n_3, A2 => l073_n_113, ZN => l073_n_170);
  l073_g12476 : ND2D1BWP7T port map(A1 => l073_n_151, A2 => l073_n_114, ZN => l073_n_168);
  l073_g12477 : INR2D1BWP7T port map(A1 => l073_n_114, B1 => l073_n_158, ZN => l073_n_167);
  l073_g12478 : AN2D1BWP7T port map(A1 => l073_n_5, A2 => l073_n_113, Z => l073_n_166);
  l073_g12479 : ND2D1BWP7T port map(A1 => l073_n_152, A2 => l073_n_114, ZN => l073_n_165);
  l073_g12480 : IND4D0BWP7T port map(A1 => l073_n_71, B1 => l073_n_72, B2 => l073_n_102, B3 => l073_n_116, ZN => l073_n_163);
  l073_g12481 : ND4D0BWP7T port map(A1 => l073_n_129, A2 => l073_n_95, A3 => l073_n_70, A4 => l073_n_60, ZN => l073_n_162);
  l073_g12482 : IND4D0BWP7T port map(A1 => l073_n_76, B1 => l073_n_77, B2 => l073_n_70, B3 => l073_n_124, ZN => l073_n_161);
  l073_g12483 : OAI222D0BWP7T port map(A1 => l073_n_145, A2 => l073_n_138, B1 => l073_n_98, B2 => l073_n_137, C1 => l073_n_104, C2 => l073_n_105, ZN => l073_n_160);
  l073_g12484 : MOAI22D0BWP7T port map(A1 => l073_n_144, A2 => l073_n_136, B1 => l073_n_138, B2 => l073_n_106, ZN => l073_n_159);
  l073_g12485 : ND3D0BWP7T port map(A1 => l073_n_140, A2 => l073_n_146, A3 => l073_n_141, ZN => l073_n_164);
  l073_g12486 : OAI211D1BWP7T port map(A1 => l073_n_13, A2 => l073_n_56, B => l073_n_143, C => l073_n_89, ZN => l073_n_157);
  l073_g12487 : INR3D0BWP7T port map(A1 => l073_n_116, B1 => l073_n_93, B2 => l073_n_125, ZN => l073_n_156);
  l073_g12488 : AOI211D1BWP7T port map(A1 => l073_n_48, A2 => y(5), B => l073_n_123, C => l073_n_109, ZN => l073_n_155);
  l073_g12489 : NR3D0BWP7T port map(A1 => l073_n_134, A2 => l073_n_46, A3 => y(4), ZN => l073_n_154);
  l073_g12490 : AO211D0BWP7T port map(A1 => l073_n_59, A2 => l073_n_11, B => l073_n_147, C => l073_n_86, Z => l073_n_153);
  l073_g12491 : ND3D0BWP7T port map(A1 => l073_n_115, A2 => l073_n_110, A3 => l073_n_45, ZN => l073_n_158);
  l073_g12494 : NR3D0BWP7T port map(A1 => l073_n_117, A2 => l073_n_45, A3 => l073_n_47, ZN => l073_n_152);
  l073_g12496 : NR3D0BWP7T port map(A1 => l073_n_122, A2 => l073_n_115, A3 => l073_n_44, ZN => l073_n_151);
  l073_g12497 : AN4D1BWP7T port map(A1 => l073_n_115, A2 => l073_n_108, A3 => l073_n_1, A4 => l073_n_45, Z => l073_n_150);
  l073_g12498 : INR2D1BWP7T port map(A1 => l073_n_118, B1 => l073_n_135, ZN => l073_n_149);
  l073_g12499 : OR2D1BWP7T port map(A1 => l073_n_134, A2 => l073_n_41, Z => l073_n_148);
  l073_g12500 : ND2D1BWP7T port map(A1 => l073_n_132, A2 => l073_n_95, ZN => l073_n_147);
  l073_g12501 : AOI211XD0BWP7T port map(A1 => l073_n_53, A2 => l073_n_33, B => l073_n_90, C => l073_n_111, ZN => l073_n_146);
  l073_g12502 : CKND1BWP7T port map(I => l073_n_144, ZN => l073_n_145);
  l073_g12503 : AOI22D0BWP7T port map(A1 => l073_n_99, A2 => y(5), B1 => l073_n_83, B2 => y_enemy3(5), ZN => l073_n_141);
  l073_g12504 : NR2XD0BWP7T port map(A1 => l073_n_123, A2 => l073_n_109, ZN => l073_n_140);
  l073_g12505 : MAOI222D1BWP7T port map(A => l073_n_88, B => x(2), C => x_enemy3(2), ZN => l073_n_144);
  l073_g12506 : NR3D0BWP7T port map(A1 => l073_n_97, A2 => l073_n_91, A3 => l073_n_69, ZN => l073_n_143);
  l073_g12507 : OAI21D0BWP7T port map(A1 => l073_n_107, A2 => l073_n_14, B => l073_n_105, ZN => l073_n_142);
  l073_g12508 : CKND1BWP7T port map(I => l073_n_136, ZN => l073_n_137);
  l073_g12509 : INVD0BWP7T port map(I => l073_n_132, ZN => l073_n_131);
  l073_g12510 : AOI211XD0BWP7T port map(A1 => l073_n_59, A2 => l073_n_25, B => l073_n_97, C => l073_n_80, ZN => l073_n_130);
  l073_g12511 : OAI21D0BWP7T port map(A1 => l073_n_74, A2 => l073_n_58, B => draw_count7(1), ZN => l073_n_129);
  l073_g12512 : AOI221D0BWP7T port map(A1 => l073_n_58, A2 => l073_n_26, B1 => l073_n_62, B2 => draw_count7(0), C => l073_n_78, ZN => l073_n_128);
  l073_g12513 : AO221D0BWP7T port map(A1 => l073_n_66, A2 => l073_n_64, B1 => l073_n_67, B2 => l073_n_27, C => l073_n_94, Z => l073_n_127);
  l073_g12514 : OA211D0BWP7T port map(A1 => l073_n_25, A2 => l073_n_60, B => l073_n_102, C => l073_n_79, Z => l073_n_126);
  l073_g12515 : OAI211D1BWP7T port map(A1 => l073_n_11, A2 => l073_n_56, B => l073_n_81, C => l073_n_75, ZN => l073_n_125);
  l073_g12516 : AOI21D0BWP7T port map(A1 => l073_n_59, A2 => l073_n_26, B => l073_n_87, ZN => l073_n_124);
  l073_g12517 : AO21D0BWP7T port map(A1 => l073_n_67, A2 => l073_n_66, B => l073_n_94, Z => l073_n_139);
  l073_g12518 : OAI22D0BWP7T port map(A1 => l073_n_68, A2 => l073_n_16, B1 => l073_n_50, B2 => x(2), ZN => l073_n_138);
  l073_g12519 : IOA21D1BWP7T port map(A1 => l073_n_50, A2 => x(2), B => l073_n_106, ZN => l073_n_136);
  l073_g12520 : ND2D1BWP7T port map(A1 => l073_n_103, A2 => l073_n_42, ZN => l073_n_135);
  l073_g12521 : ND2D1BWP7T port map(A1 => l073_n_103, A2 => l073_n_84, ZN => l073_n_134);
  l073_g12522 : IND2D1BWP7T port map(A1 => l073_n_93, B1 => l073_n_70, ZN => l073_n_133);
  l073_g12523 : INR2XD0BWP7T port map(A1 => l073_n_60, B1 => l073_n_91, ZN => l073_n_132);
  l073_g12528 : OAI22D0BWP7T port map(A1 => l073_n_52, A2 => l073_n_28, B1 => l073_n_48, B2 => y(5), ZN => l073_n_123);
  l073_g12529 : MOAI22D0BWP7T port map(A1 => l073_n_60, A2 => draw_count7(1), B1 => l073_n_74, B2 => l073_n_66, ZN => l073_n_112);
  l073_g12530 : MOAI22D0BWP7T port map(A1 => l073_n_19, A2 => y(9), B1 => l073_n_19, B2 => y(9), ZN => l073_n_111);
  l073_g12531 : MAOI22D0BWP7T port map(A1 => l073_n_84, A2 => l073_n_34, B1 => l073_n_84, B2 => l073_n_34, ZN => l073_n_122);
  l073_g12532 : MAOI22D0BWP7T port map(A1 => l073_n_43, A2 => l073_n_35, B1 => l073_n_43, B2 => l073_n_35, ZN => l073_n_121);
  l073_g12533 : MAOI22D0BWP7T port map(A1 => l073_n_43, A2 => y(3), B1 => l073_n_43, B2 => y(3), ZN => l073_n_120);
  l073_g12534 : MOAI22D0BWP7T port map(A1 => l073_n_43, A2 => l073_n_18, B1 => l073_n_43, B2 => l073_n_18, ZN => l073_n_119);
  l073_g12535 : MAOI22D0BWP7T port map(A1 => l073_n_82, A2 => y(2), B1 => l073_n_82, B2 => y(2), ZN => l073_n_118);
  l073_g12536 : ND2D1BWP7T port map(A1 => l073_n_108, A2 => l073_n_1, ZN => l073_n_110);
  l073_g12537 : MAOI22D0BWP7T port map(A1 => l073_n_42, A2 => y(1), B1 => l073_n_42, B2 => y(1), ZN => l073_n_117);
  l073_g12538 : INR3D0BWP7T port map(A1 => l073_n_79, B1 => l073_n_62, B2 => l073_n_78, ZN => l073_n_116);
  l073_g12539 : MOAI22D0BWP7T port map(A1 => l073_n_47, A2 => y(0), B1 => l073_n_47, B2 => y(0), ZN => l073_n_115);
  l073_g12540 : MAOI22D0BWP7T port map(A1 => l073_n_41, A2 => l073_n_21, B1 => l073_n_41, B2 => l073_n_21, ZN => l073_n_114);
  l073_g12541 : MOAI22D0BWP7T port map(A1 => l073_n_41, A2 => l073_n_23, B1 => l073_n_41, B2 => l073_n_23, ZN => l073_n_113);
  l073_g12542 : NR2XD0BWP7T port map(A1 => l073_n_46, A2 => l073_n_30, ZN => l073_n_101);
  l073_g12543 : NR2XD0BWP7T port map(A1 => l073_n_46, A2 => l073_n_24, ZN => l073_n_100);
  l073_g12545 : AN2D1BWP7T port map(A1 => l073_n_52, A2 => l073_n_28, Z => l073_n_109);
  l073_g12546 : ND2D1BWP7T port map(A1 => l073_n_42, A2 => l073_n_31, ZN => l073_n_108);
  l073_g12547 : NR2D0BWP7T port map(A1 => l073_n_83, A2 => y_enemy3(5), ZN => l073_n_99);
  l073_g12548 : CKAN2D1BWP7T port map(A1 => l073_n_49, A2 => l073_n_38, Z => l073_n_107);
  l073_g12549 : ND2D1BWP7T port map(A1 => l073_n_68, A2 => l073_n_16, ZN => l073_n_106);
  l073_g12550 : OR2D1BWP7T port map(A1 => l073_n_49, A2 => l073_n_15, Z => l073_n_105);
  l073_g12551 : NR2XD0BWP7T port map(A1 => l073_n_68, A2 => l073_n_16, ZN => l073_n_98);
  l073_g12552 : CKAN2D1BWP7T port map(A1 => l073_n_14, A2 => l073_n_38, Z => l073_n_104);
  l073_g12553 : INR2D1BWP7T port map(A1 => l073_n_47, B1 => l073_n_45, ZN => l073_n_103);
  l073_g12554 : NR2XD0BWP7T port map(A1 => l073_n_73, A2 => l073_n_80, ZN => l073_n_102);
  l073_g12555 : NR2D0BWP7T port map(A1 => l073_n_53, A2 => l073_n_33, ZN => l073_n_90);
  l073_g12556 : AOI22D0BWP7T port map(A1 => l073_n_59, A2 => l073_n_12, B1 => l073_n_62, B2 => l073_n_25, ZN => l073_n_89);
  l073_g12557 : AOI22D0BWP7T port map(A1 => l073_n_54, A2 => x(0), B1 => x(1), B2 => l073_n_9, ZN => l073_n_88);
  l073_g12558 : AOI21D0BWP7T port map(A1 => l073_n_57, A2 => l073_n_60, B => draw_count7(1), ZN => l073_n_87);
  l073_g12559 : OA21D0BWP7T port map(A1 => l073_n_58, A2 => l073_n_55, B => l073_n_25, Z => l073_n_86);
  l073_g12560 : AOI21D0BWP7T port map(A1 => l073_n_58, A2 => l073_n_25, B => l073_n_63, ZN => l073_n_85);
  l073_g12561 : OAI21D0BWP7T port map(A1 => l073_n_56, A2 => draw_count7(1), B => l073_n_75, ZN => l073_n_97);
  l073_g12562 : AOI21D0BWP7T port map(A1 => l073_n_62, A2 => l073_n_11, B => l073_n_59, ZN => l073_n_96);
  l073_g12563 : OAI21D0BWP7T port map(A1 => l073_n_63, A2 => l073_n_55, B => l073_n_12, ZN => l073_n_95);
  l073_g12564 : MOAI22D0BWP7T port map(A1 => l073_n_65, A2 => l073_n_26, B1 => l073_n_67, B2 => l073_n_12, ZN => l073_n_94);
  l073_g12565 : AO21D0BWP7T port map(A1 => l073_n_64, A2 => l073_n_26, B => l073_n_73, Z => l073_n_93);
  l073_g12566 : IOA21D1BWP7T port map(A1 => l073_n_58, A2 => l073_n_11, B => l073_n_77, ZN => l073_n_92);
  l073_g12567 : OAI22D0BWP7T port map(A1 => l073_n_57, A2 => l073_n_11, B1 => l073_n_60, B2 => l073_n_26, ZN => l073_n_91);
  l073_g12568 : INVD1BWP7T port map(I => l073_n_42, ZN => l073_n_84);
  l073_g12570 : INVD0BWP7T port map(I => l073_n_48, ZN => l073_n_83);
  l073_g12571 : INVD0BWP7T port map(I => l073_n_41, ZN => l073_n_82);
  l073_g12572 : ND2D1BWP7T port map(A1 => l073_n_59, A2 => draw_count7(1), ZN => l073_n_81);
  l073_g12573 : NR2D1BWP7T port map(A1 => l073_n_65, A2 => draw_count7(1), ZN => l073_n_80);
  l073_g12574 : IND2D0BWP7T port map(A1 => l073_n_13, B1 => l073_n_63, ZN => l073_n_79);
  l073_g12575 : INR2D1BWP7T port map(A1 => l073_n_59, B1 => draw_count7(1), ZN => l073_n_78);
  l073_g12576 : CKND2D0BWP7T port map(A1 => l073_n_63, A2 => l073_n_12, ZN => l073_n_77);
  l073_g12577 : NR2D0BWP7T port map(A1 => l073_n_56, A2 => l073_n_6, ZN => l073_n_76);
  l073_g12578 : NR2D0BWP7T port map(A1 => l073_n_60, A2 => l073_n_13, ZN => l073_n_69);
  l073_g12579 : CKND2D1BWP7T port map(A1 => l073_n_58, A2 => l073_n_66, ZN => l073_n_75);
  l073_g12580 : IND2D1BWP7T port map(A1 => l073_n_59, B1 => l073_n_61, ZN => l073_n_74);
  l073_g12581 : AN2D0BWP7T port map(A1 => l073_n_63, A2 => l073_n_25, Z => l073_n_73);
  l073_g12582 : ND2D1BWP7T port map(A1 => l073_n_55, A2 => l073_n_11, ZN => l073_n_72);
  l073_g12583 : INR2D1BWP7T port map(A1 => l073_n_27, B1 => l073_n_57, ZN => l073_n_71);
  l073_g12584 : ND2D1BWP7T port map(A1 => l073_n_63, A2 => l073_n_66, ZN => l073_n_70);
  l073_g12585 : INVD1BWP7T port map(I => l073_n_65, ZN => l073_n_64);
  l073_g12586 : INVD1BWP7T port map(I => l073_n_62, ZN => l073_n_61);
  l073_g12587 : INVD0BWP7T port map(I => l073_n_58, ZN => l073_n_57);
  l073_g12588 : INVD1BWP7T port map(I => l073_n_56, ZN => l073_n_55);
  l073_g12589 : IAO21D0BWP7T port map(A1 => x(1), A2 => l073_n_9, B => x_enemy3(0), ZN => l073_n_54);
  l073_g12590 : AO21D0BWP7T port map(A1 => x(4), A2 => l073_n_10, B => l073_n_14, Z => l073_n_68);
  l073_g12591 : INR2D1BWP7T port map(A1 => draw_count7(3), B1 => l073_n_32, ZN => l073_n_67);
  l073_g12592 : IND2D1BWP7T port map(A1 => l073_n_27, B1 => l073_n_13, ZN => l073_n_66);
  l073_g12593 : ND2D1BWP7T port map(A1 => l073_n_39, A2 => draw_count7(3), ZN => l073_n_65);
  l073_g12594 : NR2D1BWP7T port map(A1 => l073_n_32, A2 => draw_count7(3), ZN => l073_n_63);
  l073_g12595 : INR2D1BWP7T port map(A1 => l073_n_22, B1 => draw_count7(3), ZN => l073_n_62);
  l073_g12596 : ND2D1BWP7T port map(A1 => l073_n_36, A2 => draw_count7(3), ZN => l073_n_60);
  l073_g12597 : NR2D1BWP7T port map(A1 => l073_n_37, A2 => draw_count7(3), ZN => l073_n_59);
  l073_g12598 : NR2D1BWP7T port map(A1 => l073_n_40, A2 => draw_count7(3), ZN => l073_n_58);
  l073_g12599 : ND2D1BWP7T port map(A1 => l073_n_22, A2 => draw_count7(3), ZN => l073_n_56);
  l073_g12601 : INVD0BWP7T port map(I => l073_n_45, ZN => l073_n_44);
  l073_g12602 : MOAI22D0BWP7T port map(A1 => y(8), A2 => y_enemy3(8), B1 => y(8), B2 => y_enemy3(8), ZN => l073_n_53);
  l073_g12603 : MAOI22D0BWP7T port map(A1 => y(7), A2 => y_enemy3(7), B1 => y(7), B2 => y_enemy3(7), ZN => l073_n_52);
  l073_g12604 : MOAI22D0BWP7T port map(A1 => x(7), A2 => x_enemy3(7), B1 => x(7), B2 => x_enemy3(7), ZN => l073_n_51);
  l073_g12605 : MAOI22D0BWP7T port map(A1 => x(3), A2 => x_enemy3(3), B1 => x(3), B2 => x_enemy3(3), ZN => l073_n_50);
  l073_g12606 : MAOI22D0BWP7T port map(A1 => x(6), A2 => x_enemy3(6), B1 => x(6), B2 => x_enemy3(6), ZN => l073_n_49);
  l073_g12607 : OAI21D0BWP7T port map(A1 => l073_n_7, A2 => y_enemy3(6), B => l073_n_28, ZN => l073_n_48);
  l073_g12608 : MOAI22D0BWP7T port map(A1 => y(1), A2 => y_enemy3(1), B1 => y(1), B2 => y_enemy3(1), ZN => l073_n_47);
  l073_g12609 : MAOI22D0BWP7T port map(A1 => y(5), A2 => y_enemy3(5), B1 => y(5), B2 => y_enemy3(5), ZN => l073_n_46);
  l073_g12610 : MAOI22D0BWP7T port map(A1 => y(0), A2 => y_enemy3(0), B1 => y(0), B2 => y_enemy3(0), ZN => l073_n_45);
  l073_g12611 : MOAI22D0BWP7T port map(A1 => y(4), A2 => y_enemy3(4), B1 => y(4), B2 => y_enemy3(4), ZN => l073_n_43);
  l073_g12612 : MAOI22D0BWP7T port map(A1 => y(2), A2 => y_enemy3(2), B1 => y(2), B2 => y_enemy3(2), ZN => l073_n_42);
  l073_g12613 : MOAI22D0BWP7T port map(A1 => y(3), A2 => y_enemy3(3), B1 => y(3), B2 => y_enemy3(3), ZN => l073_n_41);
  l073_g12614 : INVD0BWP7T port map(I => l073_n_39, ZN => l073_n_40);
  l073_g12615 : CKND1BWP7T port map(I => l073_n_36, ZN => l073_n_37);
  l073_g12616 : INVD1BWP7T port map(I => l073_n_26, ZN => l073_n_25);
  l073_g12617 : INR2D1BWP7T port map(A1 => draw_count7(4), B1 => draw_count7(2), ZN => l073_n_39);
  l073_g12618 : IND2D1BWP7T port map(A1 => x_enemy3(5), B1 => x(5), ZN => l073_n_38);
  l073_g12619 : INR2D1BWP7T port map(A1 => draw_count7(2), B1 => draw_count7(4), ZN => l073_n_36);
  l073_g12620 : IND2D0BWP7T port map(A1 => y_enemy3(3), B1 => y(3), ZN => l073_n_35);
  l073_g12621 : IND2D1BWP7T port map(A1 => y_enemy3(1), B1 => y(1), ZN => l073_n_34);
  l073_g12622 : INR2XD0BWP7T port map(A1 => y_enemy3(7), B1 => y(7), ZN => l073_n_33);
  l073_g12623 : ND2D1BWP7T port map(A1 => draw_count7(2), A2 => draw_count7(4), ZN => l073_n_32);
  l073_g12624 : IND2D1BWP7T port map(A1 => y(1), B1 => y_enemy3(1), ZN => l073_n_31);
  l073_g12625 : IND2D1BWP7T port map(A1 => y_enemy3(4), B1 => y(4), ZN => l073_n_30);
  l073_g12626 : IND2D1BWP7T port map(A1 => x(7), B1 => x_enemy3(7), ZN => l073_n_29);
  l073_g12627 : ND2D1BWP7T port map(A1 => l073_n_7, A2 => y_enemy3(6), ZN => l073_n_28);
  l073_g12628 : INR2D1BWP7T port map(A1 => draw_count7(0), B1 => draw_count7(1), ZN => l073_n_27);
  l073_g12629 : CKND2D1BWP7T port map(A1 => draw_count7(1), A2 => draw_count7(0), ZN => l073_n_26);
  l073_g12630 : INVD1BWP7T port map(I => l073_n_12, ZN => l073_n_11);
  l073_g12631 : INR2D1BWP7T port map(A1 => y_enemy3(4), B1 => y(4), ZN => l073_n_24);
  l073_g12632 : IND2D1BWP7T port map(A1 => y(2), B1 => y_enemy3(2), ZN => l073_n_23);
  l073_g12633 : NR2D0BWP7T port map(A1 => draw_count7(2), A2 => draw_count7(4), ZN => l073_n_22);
  l073_g12634 : IND2D1BWP7T port map(A1 => y_enemy3(2), B1 => y(2), ZN => l073_n_21);
  l073_g12635 : NR2D0BWP7T port map(A1 => l073_n_8, A2 => x_enemy3(8), ZN => l073_n_20);
  l073_g12636 : IND2D1BWP7T port map(A1 => y(8), B1 => y_enemy3(8), ZN => l073_n_19);
  l073_g12637 : IND2D1BWP7T port map(A1 => y(3), B1 => y_enemy3(3), ZN => l073_n_18);
  l073_g12638 : IND2D1BWP7T port map(A1 => x_enemy3(6), B1 => x(6), ZN => l073_n_17);
  l073_g12639 : IND2D1BWP7T port map(A1 => x(3), B1 => x_enemy3(3), ZN => l073_n_16);
  l073_g12640 : INR2XD0BWP7T port map(A1 => x_enemy3(5), B1 => x(5), ZN => l073_n_15);
  l073_g12641 : NR2D0BWP7T port map(A1 => x(4), A2 => l073_n_10, ZN => l073_n_14);
  l073_g12642 : IND2D1BWP7T port map(A1 => draw_count7(0), B1 => draw_count7(1), ZN => l073_n_13);
  l073_g12643 : NR2D0BWP7T port map(A1 => draw_count7(1), A2 => draw_count7(0), ZN => l073_n_12);
  l073_g12644 : CKND1BWP7T port map(I => x_enemy3(4), ZN => l073_n_10);
  l073_g12645 : INVD0BWP7T port map(I => x_enemy3(1), ZN => l073_n_9);
  l073_g12646 : CKND1BWP7T port map(I => x(8), ZN => l073_n_8);
  l073_g12647 : CKND1BWP7T port map(I => y(6), ZN => l073_n_7);
  l073_g12648 : INVD0BWP7T port map(I => draw_count7(1), ZN => l073_n_6);
  l073_g2 : INR3D0BWP7T port map(A1 => l073_n_122, B1 => l073_n_115, B2 => l073_n_44, ZN => l073_n_5);
  l073_g12649 : IND2D1BWP7T port map(A1 => l073_n_119, B1 => l073_n_177, ZN => l073_n_4);
  l073_g12650 : INR3D0BWP7T port map(A1 => l073_n_117, B1 => l073_n_45, B2 => l073_n_47, ZN => l073_n_3);
  l073_g12651 : IIND4D0BWP7T port map(A1 => l073_n_121, A2 => l073_n_113, B1 => l073_n_150, B2 => l073_n_177, ZN => l073_n_2);
  l073_g12652 : IND2D1BWP7T port map(A1 => l073_n_31, B1 => l073_n_84, ZN => l073_n_1);
  l073_g12653 : INR3D0BWP7T port map(A1 => l073_n_46, B1 => l073_n_134, B2 => l073_n_82, ZN => l073_n_0);
  l02_count_reg_9 : DFQD1BWP7T port map(CP => clk, D => l02_n_39, Q => y(9));
  l02_g1019 : AO22D0BWP7T port map(A1 => l02_n_1, A2 => y(9), B1 => l02_n_22, B2 => l02_n_37, Z => l02_n_39);
  l02_g1020 : AO21D0BWP7T port map(A1 => l02_n_1, A2 => y(8), B => l02_n_36, Z => l02_n_38);
  l02_count_reg_7 : DFQD1BWP7T port map(CP => clk, D => l02_n_35, Q => y(7));
  l02_g1022 : OAI31D0BWP7T port map(A1 => y(9), A2 => l02_n_5, A3 => l02_n_31, B => l02_n_6, ZN => l02_n_37);
  l02_g1023 : NR3D0BWP7T port map(A1 => l02_n_21, A2 => l02_n_31, A3 => y(8), ZN => l02_n_36);
  l02_g1024 : MOAI22D0BWP7T port map(A1 => l02_n_21, A2 => l02_n_32, B1 => l02_n_14, B2 => y(7), ZN => l02_n_35);
  l02_g1028 : OAI22D0BWP7T port map(A1 => l02_n_29, A2 => l02_n_3, B1 => l02_n_21, B2 => l02_n_30, ZN => l02_n_34);
  l02_g1029 : OAI32D1BWP7T port map(A1 => y(5), A2 => l02_n_19, A3 => l02_n_21, B1 => l02_n_4, B2 => l02_n_29, ZN => l02_n_33);
  l02_g1030 : MAOI22D0BWP7T port map(A1 => l02_n_28, A2 => y(7), B1 => l02_n_28, B2 => y(7), ZN => l02_n_32);
  l02_count_reg_4 : DFQD1BWP7T port map(CP => clk, D => l02_n_27, Q => y(4));
  l02_g1032 : MAOI22D0BWP7T port map(A1 => l02_n_4, A2 => y(6), B1 => l02_n_26, B2 => y(6), ZN => l02_n_30);
  l02_g1033 : IND2D1BWP7T port map(A1 => l02_n_28, B1 => y(7), ZN => l02_n_31);
  l02_count_reg_1 : DFQD1BWP7T port map(CP => clk, D => l02_n_25, Q => y(1));
  l02_count_reg_3 : DFQD1BWP7T port map(CP => clk, D => l02_n_23, Q => y(3));
  l02_count_reg_2 : DFQD1BWP7T port map(CP => clk, D => l02_n_24, Q => y(2));
  l02_g1037 : MOAI22D0BWP7T port map(A1 => l02_n_21, A2 => l02_n_20, B1 => l02_n_14, B2 => y(4), ZN => l02_n_27);
  l02_g1038 : AOI21D0BWP7T port map(A1 => l02_n_22, A2 => l02_n_19, B => l02_n_14, ZN => l02_n_29);
  l02_g1039 : OR2D1BWP7T port map(A1 => l02_n_26, A2 => l02_n_3, Z => l02_n_28);
  l02_count_reg_0 : DFXQD1BWP7T port map(CP => clk, DA => l02_n_14, DB => l02_n_22, SA => y(0), Q => y(0));
  l02_g1041 : MOAI22D0BWP7T port map(A1 => l02_n_21, A2 => l02_n_0, B1 => l02_n_14, B2 => y(1), ZN => l02_n_25);
  l02_g1042 : OR2D1BWP7T port map(A1 => l02_n_19, A2 => l02_n_4, Z => l02_n_26);
  l02_g1043 : MOAI22D0BWP7T port map(A1 => l02_n_21, A2 => l02_n_13, B1 => l02_n_14, B2 => y(2), ZN => l02_n_24);
  l02_g1044 : MOAI22D0BWP7T port map(A1 => l02_n_21, A2 => l02_n_17, B1 => l02_n_14, B2 => y(3), ZN => l02_n_23);
  l02_g1045 : INVD1BWP7T port map(I => l02_n_22, ZN => l02_n_21);
  l02_g1046 : NR3D0BWP7T port map(A1 => l02_n_18, A2 => l02_n_11, A3 => reset, ZN => l02_n_22);
  l02_g1047 : MAOI22D0BWP7T port map(A1 => l02_n_16, A2 => y(4), B1 => l02_n_16, B2 => y(4), ZN => l02_n_20);
  l02_g1048 : IND2D1BWP7T port map(A1 => l02_n_16, B1 => y(4), ZN => l02_n_19);
  l02_g1049 : NR4D0BWP7T port map(A1 => l02_n_15, A2 => y(7), A3 => y(6), A4 => y(5), ZN => l02_n_18);
  l02_g1050 : MAOI22D0BWP7T port map(A1 => l02_n_12, A2 => y(3), B1 => l02_n_12, B2 => y(3), ZN => l02_n_17);
  l02_g1051 : IND2D1BWP7T port map(A1 => l02_n_12, B1 => y(3), ZN => l02_n_16);
  l02_g1052 : IND4D0BWP7T port map(A1 => y(4), B1 => y(2), B2 => y(3), B3 => l02_n_10, ZN => l02_n_15);
  l02_g1054 : INR2XD0BWP7T port map(A1 => l02_n_11, B1 => reset, ZN => l02_n_14);
  l02_g1055 : MAOI22D0BWP7T port map(A1 => l02_n_7, A2 => y(2), B1 => l02_n_7, B2 => y(2), ZN => l02_n_13);
  l02_g1056 : IND2D1BWP7T port map(A1 => l02_n_7, B1 => y(2), ZN => l02_n_12);
  l02_g1057 : IND4D0BWP7T port map(A1 => l02_n_9, B1 => x(1), B2 => x(2), B3 => l02_n_8, ZN => l02_n_11);
  l02_g1058 : NR3D0BWP7T port map(A1 => l02_n_6, A2 => y(1), A3 => y(0), ZN => l02_n_10);
  l02_g1059 : ND3D0BWP7T port map(A1 => x(8), A2 => x(7), A3 => x(0), ZN => l02_n_9);
  l02_g1060 : INR4D0BWP7T port map(A1 => x(3), B1 => x(6), B2 => x(4), B3 => x(5), ZN => l02_n_8);
  l02_g1062 : ND2D1BWP7T port map(A1 => y(1), A2 => y(0), ZN => l02_n_7);
  l02_g1063 : ND2D1BWP7T port map(A1 => l02_n_5, A2 => y(9), ZN => l02_n_6);
  l02_g2 : AO21D0BWP7T port map(A1 => l02_n_22, A2 => l02_n_31, B => l02_n_14, Z => l02_n_1);
  l02_g1074 : XNR2D1BWP7T port map(A1 => y(1), A2 => y(0), ZN => l02_n_0);
  l02_count_reg_8 : DFD1BWP7T port map(CP => clk, D => l02_n_38, Q => y(8), QN => l02_n_5);
  l02_count_reg_5 : DFD1BWP7T port map(CP => clk, D => l02_n_33, Q => y(5), QN => l02_n_4);
  l02_count_reg_6 : DFD1BWP7T port map(CP => clk, D => l02_n_34, Q => y(6), QN => l02_n_3);
  l074_g12411 : OAI221D0BWP7T port map(A1 => l074_n_221, A2 => l074_n_183, B1 => l074_n_155, B2 => l074_n_224, C => l074_n_245, ZN => r8);
  l074_g12412 : NR4D0BWP7T port map(A1 => l074_n_244, A2 => l074_n_234, A3 => l074_n_228, A4 => l074_n_205, ZN => l074_n_245);
  l074_g12413 : IND4D0BWP7T port map(A1 => l074_n_232, B1 => l074_n_227, B2 => l074_n_233, B3 => l074_n_241, ZN => l074_n_244);
  l074_g12414 : AO211D0BWP7T port map(A1 => l074_n_217, A2 => l074_n_91, B => l074_n_242, C => l074_n_240, Z => g8);
  l074_g12415 : OAI211D1BWP7T port map(A1 => l074_n_125, A2 => l074_n_221, B => l074_n_238, C => l074_n_230, ZN => l074_n_242);
  l074_g12416 : MAOI22D0BWP7T port map(A1 => l074_n_214, A2 => l074_n_161, B1 => l074_n_235, B2 => l074_n_193, ZN => l074_n_241);
  l074_g12417 : AO221D0BWP7T port map(A1 => l074_n_214, A2 => l074_n_138, B1 => l074_n_211, B2 => l074_n_126, C => l074_n_236, Z => l074_n_240);
  l074_g12418 : OAI32D1BWP7T port map(A1 => l074_n_26, A2 => l074_n_61, A3 => l074_n_221, B1 => l074_n_95, B2 => l074_n_223, ZN => b8);
  l074_g12419 : AOI211XD0BWP7T port map(A1 => l074_n_198, A2 => l074_n_70, B => l074_n_231, C => l074_n_225, ZN => l074_n_238);
  l074_g12420 : ND3D0BWP7T port map(A1 => l074_n_219, A2 => l074_n_210, A3 => l074_n_197, ZN => enable8);
  l074_g12421 : OAI211D1BWP7T port map(A1 => l074_n_84, A2 => l074_n_203, B => l074_n_218, C => l074_n_226, ZN => l074_n_236);
  l074_g12422 : ND4D0BWP7T port map(A1 => l074_n_215, A2 => l074_n_186, A3 => l074_n_180, A4 => l074_n_164, ZN => l074_n_235);
  l074_g12423 : OAI211D1BWP7T port map(A1 => l074_n_171, A2 => l074_n_223, B => l074_n_220, C => l074_n_206, ZN => l074_n_234);
  l074_g12424 : AOI22D0BWP7T port map(A1 => l074_n_211, A2 => l074_n_156, B1 => l074_n_216, B2 => l074_n_160, ZN => l074_n_233);
  l074_g12425 : AOI31D0BWP7T port map(A1 => l074_n_129, A2 => l074_n_131, A3 => l074_n_61, B => l074_n_229, ZN => l074_n_232);
  l074_g12426 : AOI21D0BWP7T port map(A1 => l074_n_131, A2 => l074_n_71, B => l074_n_224, ZN => l074_n_231);
  l074_g12427 : OAI21D0BWP7T port map(A1 => l074_n_132, A2 => l074_n_91, B => l074_n_222, ZN => l074_n_230);
  l074_g12428 : AOI21D0BWP7T port map(A1 => l074_n_209, A2 => l074_n_149, B => l074_n_195, ZN => l074_n_229);
  l074_g12429 : IAO21D0BWP7T port map(A1 => l074_n_152, A2 => l074_n_70, B => l074_n_212, ZN => l074_n_228);
  l074_g12430 : OAI31D0BWP7T port map(A1 => l074_n_75, A2 => l074_n_91, A3 => l074_n_111, B => l074_n_213, ZN => l074_n_227);
  l074_g12431 : OAI21D0BWP7T port map(A1 => l074_n_132, A2 => l074_n_138, B => l074_n_213, ZN => l074_n_226);
  l074_g12432 : AOI21D0BWP7T port map(A1 => l074_n_101, A2 => l074_n_69, B => l074_n_212, ZN => l074_n_225);
  l074_g12433 : INVD0BWP7T port map(I => l074_n_222, ZN => l074_n_223);
  l074_g12434 : OAI21D0BWP7T port map(A1 => l074_n_90, A2 => l074_n_55, B => l074_n_217, ZN => l074_n_220);
  l074_g12435 : AOI22D0BWP7T port map(A1 => l074_n_204, A2 => l074_n_192, B1 => l074_n_202, B2 => l074_n_177, ZN => l074_n_219);
  l074_g12436 : OAI21D0BWP7T port map(A1 => l074_n_92, A2 => l074_n_64, B => l074_n_216, ZN => l074_n_218);
  l074_g12437 : AOI22D0BWP7T port map(A1 => l074_n_208, A2 => l074_n_150, B1 => l074_n_209, B2 => l074_n_4, ZN => l074_n_224);
  l074_g12438 : OAI32D1BWP7T port map(A1 => l074_n_117, A2 => l074_n_134, A3 => l074_n_197, B1 => l074_n_157, B2 => l074_n_207, ZN => l074_n_222);
  l074_g12439 : AOI22D0BWP7T port map(A1 => l074_n_209, A2 => l074_n_6, B1 => l074_n_208, B2 => l074_n_151, ZN => l074_n_221);
  l074_g12440 : AOI211D1BWP7T port map(A1 => l074_n_127, A2 => l074_n_56, B => l074_n_196, C => l074_n_187, ZN => l074_n_215);
  l074_g12441 : OAI22D0BWP7T port map(A1 => l074_n_199, A2 => l074_n_170, B1 => l074_n_193, B2 => l074_n_180, ZN => l074_n_217);
  l074_g12442 : IOA21D1BWP7T port map(A1 => l074_n_202, A2 => l074_n_166, B => l074_n_210, ZN => l074_n_216);
  l074_g12443 : MOAI22D0BWP7T port map(A1 => l074_n_199, A2 => l074_n_164, B1 => l074_n_202, B2 => l074_n_165, ZN => l074_n_214);
  l074_g12444 : MOAI22D0BWP7T port map(A1 => l074_n_199, A2 => l074_n_167, B1 => l074_n_202, B2 => l074_n_168, ZN => l074_n_213);
  l074_g12445 : MAOI22D0BWP7T port map(A1 => l074_n_200, A2 => l074_n_165, B1 => l074_n_201, B2 => l074_n_164, ZN => l074_n_212);
  l074_g12446 : MOAI22D0BWP7T port map(A1 => l074_n_193, A2 => l074_n_186, B1 => l074_n_200, B2 => l074_n_166, ZN => l074_n_211);
  l074_g12447 : INVD0BWP7T port map(I => l074_n_208, ZN => l074_n_207);
  l074_g12448 : ND2D1BWP7T port map(A1 => l074_n_200, A2 => l074_n_148, ZN => l074_n_210);
  l074_g12449 : NR2D1BWP7T port map(A1 => l074_n_197, A2 => l074_n_112, ZN => l074_n_209);
  l074_g12450 : NR2D1BWP7T port map(A1 => l074_n_197, A2 => l074_n_113, ZN => l074_n_208);
  l074_g12451 : OAI21D0BWP7T port map(A1 => l074_n_130, A2 => l074_n_75, B => l074_n_198, ZN => l074_n_206);
  l074_g12452 : AOI21D0BWP7T port map(A1 => l074_n_142, A2 => l074_n_80, B => l074_n_203, ZN => l074_n_205);
  l074_g12453 : ND4D0BWP7T port map(A1 => l074_n_194, A2 => l074_n_189, A3 => l074_n_3, A4 => l074_n_181, ZN => l074_n_204);
  l074_g12454 : INVD0BWP7T port map(I => l074_n_202, ZN => l074_n_201);
  l074_g12455 : INVD0BWP7T port map(I => l074_n_200, ZN => l074_n_199);
  l074_g12456 : CKND2D1BWP7T port map(A1 => l074_n_192, A2 => l074_n_187, ZN => l074_n_203);
  l074_g12457 : NR2D1BWP7T port map(A1 => l074_n_193, A2 => l074_n_184, ZN => l074_n_202);
  l074_g12458 : NR2D1BWP7T port map(A1 => l074_n_193, A2 => l074_n_5, ZN => l074_n_200);
  l074_g12459 : OA31D1BWP7T port map(A1 => l074_n_119, A2 => l074_n_147, A3 => l074_n_174, B => l074_n_194, Z => l074_n_196);
  l074_g12460 : NR4D0BWP7T port map(A1 => l074_n_193, A2 => l074_n_172, A3 => l074_n_163, A4 => l074_n_43, ZN => l074_n_195);
  l074_g12461 : AOI21D0BWP7T port map(A1 => l074_n_3, A2 => l074_n_181, B => l074_n_193, ZN => l074_n_198);
  l074_g12462 : ND3D0BWP7T port map(A1 => l074_n_192, A2 => l074_n_175, A3 => l074_n_120, ZN => l074_n_197);
  l074_g12463 : INR2XD0BWP7T port map(A1 => l074_n_186, B1 => l074_n_191, ZN => l074_n_194);
  l074_g12464 : INVD1BWP7T port map(I => l074_n_193, ZN => l074_n_192);
  l074_g12465 : OAI221D0BWP7T port map(A1 => l074_n_173, A2 => l074_n_141, B1 => l074_n_30, B2 => l074_n_21, C => l074_n_190, ZN => l074_n_193);
  l074_g12466 : OAI221D0BWP7T port map(A1 => l074_n_5, A2 => l074_n_178, B1 => l074_n_170, B2 => l074_n_184, C => l074_n_180, ZN => l074_n_191);
  l074_g12467 : AOI221D0BWP7T port map(A1 => l074_n_9, A2 => x_enemy4(8), B1 => l074_n_51, B2 => l074_n_18, C => l074_n_185, ZN => l074_n_190);
  l074_g12468 : IAO21D0BWP7T port map(A1 => l074_n_184, A2 => l074_n_182, B => l074_n_188, ZN => l074_n_189);
  l074_g12469 : AOI21D0BWP7T port map(A1 => l074_n_182, A2 => l074_n_170, B => l074_n_5, ZN => l074_n_188);
  l074_g12470 : OAI22D0BWP7T port map(A1 => l074_n_184, A2 => l074_n_167, B1 => l074_n_5, B2 => l074_n_169, ZN => l074_n_187);
  l074_g12471 : IND2D1BWP7T port map(A1 => l074_n_184, B1 => l074_n_148, ZN => l074_n_186);
  l074_g12472 : AO21D0BWP7T port map(A1 => l074_n_21, A2 => l074_n_30, B => l074_n_179, Z => l074_n_185);
  l074_g12474 : NR3D0BWP7T port map(A1 => l074_n_162, A2 => l074_n_90, A3 => l074_n_64, ZN => l074_n_183);
  l074_g12476 : ND2D1BWP7T port map(A1 => l074_n_176, A2 => l074_n_118, ZN => l074_n_184);
  l074_g12477 : MOAI22D0BWP7T port map(A1 => l074_n_51, A2 => l074_n_18, B1 => l074_n_159, B2 => l074_n_141, ZN => l074_n_179);
  l074_g12478 : INR3D0BWP7T port map(A1 => l074_n_167, B1 => l074_n_165, B2 => l074_n_166, ZN => l074_n_182);
  l074_g12479 : ND4D0BWP7T port map(A1 => l074_n_1, A2 => l074_n_154, A3 => l074_n_145, A4 => l074_n_43, ZN => l074_n_181);
  l074_g12480 : IND3D1BWP7T port map(A1 => l074_n_147, B1 => l074_n_119, B2 => l074_n_176, ZN => l074_n_180);
  l074_g12481 : CKND1BWP7T port map(I => l074_n_177, ZN => l074_n_178);
  l074_g12482 : INVD0BWP7T port map(I => l074_n_175, ZN => l074_n_174);
  l074_g12483 : ND2D1BWP7T port map(A1 => l074_n_169, A2 => l074_n_164, ZN => l074_n_177);
  l074_g12484 : AOI211XD0BWP7T port map(A1 => l074_n_46, A2 => l074_n_31, B => l074_n_163, C => l074_n_100, ZN => l074_n_176);
  l074_g12485 : AOI211XD0BWP7T port map(A1 => l074_n_46, A2 => l074_n_25, B => l074_n_163, C => l074_n_99, ZN => l074_n_175);
  l074_g12486 : AOI221D0BWP7T port map(A1 => l074_n_106, A2 => l074_n_16, B1 => l074_n_49, B2 => l074_n_103, C => l074_n_158, ZN => l074_n_173);
  l074_g12487 : AOI22D0BWP7T port map(A1 => l074_n_1, A2 => y(4), B1 => l074_n_153, B2 => l074_n_41, ZN => l074_n_172);
  l074_g12488 : INR4D0BWP7T port map(A1 => l074_n_95, B1 => l074_n_93, B2 => l074_n_146, B3 => l074_n_132, ZN => l074_n_171);
  l074_g12489 : INVD0BWP7T port map(I => l074_n_169, ZN => l074_n_168);
  l074_g12490 : ND2D1BWP7T port map(A1 => l074_n_149, A2 => l074_n_112, ZN => l074_n_170);
  l074_g12491 : ND2D1BWP7T port map(A1 => l074_n_4, A2 => l074_n_112, ZN => l074_n_169);
  l074_g12492 : ND2D1BWP7T port map(A1 => l074_n_150, A2 => l074_n_113, ZN => l074_n_167);
  l074_g12493 : INR2D1BWP7T port map(A1 => l074_n_113, B1 => l074_n_157, ZN => l074_n_166);
  l074_g12494 : AN2D1BWP7T port map(A1 => l074_n_6, A2 => l074_n_112, Z => l074_n_165);
  l074_g12495 : ND2D1BWP7T port map(A1 => l074_n_151, A2 => l074_n_113, ZN => l074_n_164);
  l074_g12496 : IND4D0BWP7T port map(A1 => l074_n_70, B1 => l074_n_71, B2 => l074_n_101, B3 => l074_n_115, ZN => l074_n_162);
  l074_g12497 : ND4D0BWP7T port map(A1 => l074_n_128, A2 => l074_n_94, A3 => l074_n_69, A4 => l074_n_60, ZN => l074_n_161);
  l074_g12498 : IND4D0BWP7T port map(A1 => l074_n_75, B1 => l074_n_69, B2 => l074_n_76, B3 => l074_n_123, ZN => l074_n_160);
  l074_g12499 : OAI222D0BWP7T port map(A1 => l074_n_144, A2 => l074_n_137, B1 => l074_n_97, B2 => l074_n_136, C1 => l074_n_103, C2 => l074_n_104, ZN => l074_n_159);
  l074_g12500 : MOAI22D0BWP7T port map(A1 => l074_n_143, A2 => l074_n_135, B1 => l074_n_137, B2 => l074_n_105, ZN => l074_n_158);
  l074_g12501 : ND3D0BWP7T port map(A1 => l074_n_139, A2 => l074_n_145, A3 => l074_n_140, ZN => l074_n_163);
  l074_g12502 : OAI211D1BWP7T port map(A1 => l074_n_14, A2 => l074_n_56, B => l074_n_142, C => l074_n_88, ZN => l074_n_156);
  l074_g12503 : INR3D0BWP7T port map(A1 => l074_n_115, B1 => l074_n_92, B2 => l074_n_124, ZN => l074_n_155);
  l074_g12504 : AOI211D1BWP7T port map(A1 => l074_n_48, A2 => y(5), B => l074_n_122, C => l074_n_108, ZN => l074_n_154);
  l074_g12505 : NR3D0BWP7T port map(A1 => l074_n_133, A2 => l074_n_46, A3 => y(4), ZN => l074_n_153);
  l074_g12506 : AO211D0BWP7T port map(A1 => l074_n_59, A2 => l074_n_12, B => l074_n_146, C => l074_n_85, Z => l074_n_152);
  l074_g12507 : ND3D0BWP7T port map(A1 => l074_n_114, A2 => l074_n_109, A3 => l074_n_45, ZN => l074_n_157);
  l074_g12510 : NR3D0BWP7T port map(A1 => l074_n_116, A2 => l074_n_45, A3 => l074_n_47, ZN => l074_n_151);
  l074_g12512 : NR3D0BWP7T port map(A1 => l074_n_121, A2 => l074_n_114, A3 => l074_n_44, ZN => l074_n_150);
  l074_g12513 : AN4D1BWP7T port map(A1 => l074_n_114, A2 => l074_n_107, A3 => l074_n_2, A4 => l074_n_45, Z => l074_n_149);
  l074_g12514 : INR2D1BWP7T port map(A1 => l074_n_117, B1 => l074_n_134, ZN => l074_n_148);
  l074_g12515 : OR2D1BWP7T port map(A1 => l074_n_133, A2 => l074_n_41, Z => l074_n_147);
  l074_g12516 : ND2D1BWP7T port map(A1 => l074_n_131, A2 => l074_n_94, ZN => l074_n_146);
  l074_g12517 : AOI211XD0BWP7T port map(A1 => l074_n_53, A2 => l074_n_34, B => l074_n_89, C => l074_n_110, ZN => l074_n_145);
  l074_g12518 : CKND1BWP7T port map(I => l074_n_143, ZN => l074_n_144);
  l074_g12519 : AOI22D0BWP7T port map(A1 => l074_n_98, A2 => y(5), B1 => l074_n_82, B2 => y_enemy4(5), ZN => l074_n_140);
  l074_g12520 : NR2XD0BWP7T port map(A1 => l074_n_122, A2 => l074_n_108, ZN => l074_n_139);
  l074_g12521 : MAOI222D1BWP7T port map(A => l074_n_87, B => x(2), C => x_enemy4(2), ZN => l074_n_143);
  l074_g12522 : NR3D0BWP7T port map(A1 => l074_n_96, A2 => l074_n_90, A3 => l074_n_68, ZN => l074_n_142);
  l074_g12523 : OAI21D0BWP7T port map(A1 => l074_n_106, A2 => l074_n_15, B => l074_n_104, ZN => l074_n_141);
  l074_g12524 : CKND1BWP7T port map(I => l074_n_135, ZN => l074_n_136);
  l074_g12525 : INVD0BWP7T port map(I => l074_n_131, ZN => l074_n_130);
  l074_g12526 : AOI211XD0BWP7T port map(A1 => l074_n_59, A2 => l074_n_26, B => l074_n_96, C => l074_n_79, ZN => l074_n_129);
  l074_g12527 : OAI21D0BWP7T port map(A1 => l074_n_73, A2 => l074_n_58, B => draw_count8(1), ZN => l074_n_128);
  l074_g12528 : AOI221D0BWP7T port map(A1 => l074_n_58, A2 => l074_n_27, B1 => l074_n_62, B2 => draw_count8(0), C => l074_n_77, ZN => l074_n_127);
  l074_g12529 : AO221D0BWP7T port map(A1 => l074_n_65, A2 => l074_n_64, B1 => l074_n_66, B2 => l074_n_28, C => l074_n_93, Z => l074_n_126);
  l074_g12530 : OA211D0BWP7T port map(A1 => l074_n_26, A2 => l074_n_60, B => l074_n_101, C => l074_n_78, Z => l074_n_125);
  l074_g12531 : OAI211D1BWP7T port map(A1 => l074_n_12, A2 => l074_n_56, B => l074_n_80, C => l074_n_74, ZN => l074_n_124);
  l074_g12532 : AOI21D0BWP7T port map(A1 => l074_n_59, A2 => l074_n_27, B => l074_n_86, ZN => l074_n_123);
  l074_g12533 : AO21D0BWP7T port map(A1 => l074_n_66, A2 => l074_n_65, B => l074_n_93, Z => l074_n_138);
  l074_g12534 : OAI22D0BWP7T port map(A1 => l074_n_67, A2 => l074_n_17, B1 => l074_n_50, B2 => x(2), ZN => l074_n_137);
  l074_g12535 : IOA21D1BWP7T port map(A1 => l074_n_50, A2 => x(2), B => l074_n_105, ZN => l074_n_135);
  l074_g12536 : ND2D1BWP7T port map(A1 => l074_n_102, A2 => l074_n_42, ZN => l074_n_134);
  l074_g12537 : ND2D1BWP7T port map(A1 => l074_n_102, A2 => l074_n_83, ZN => l074_n_133);
  l074_g12538 : IND2D1BWP7T port map(A1 => l074_n_92, B1 => l074_n_69, ZN => l074_n_132);
  l074_g12539 : INR2XD0BWP7T port map(A1 => l074_n_60, B1 => l074_n_90, ZN => l074_n_131);
  l074_g12544 : OAI22D0BWP7T port map(A1 => l074_n_52, A2 => l074_n_29, B1 => l074_n_48, B2 => y(5), ZN => l074_n_122);
  l074_g12545 : MOAI22D0BWP7T port map(A1 => l074_n_60, A2 => draw_count8(1), B1 => l074_n_73, B2 => l074_n_65, ZN => l074_n_111);
  l074_g12546 : MOAI22D0BWP7T port map(A1 => l074_n_20, A2 => y(9), B1 => l074_n_20, B2 => y(9), ZN => l074_n_110);
  l074_g12547 : MAOI22D0BWP7T port map(A1 => l074_n_83, A2 => l074_n_35, B1 => l074_n_83, B2 => l074_n_35, ZN => l074_n_121);
  l074_g12548 : MAOI22D0BWP7T port map(A1 => l074_n_43, A2 => l074_n_36, B1 => l074_n_43, B2 => l074_n_36, ZN => l074_n_120);
  l074_g12549 : MAOI22D0BWP7T port map(A1 => l074_n_43, A2 => y(3), B1 => l074_n_43, B2 => y(3), ZN => l074_n_119);
  l074_g12550 : MAOI22D0BWP7T port map(A1 => l074_n_43, A2 => l074_n_19, B1 => l074_n_43, B2 => l074_n_19, ZN => l074_n_118);
  l074_g12551 : MAOI22D0BWP7T port map(A1 => l074_n_81, A2 => y(2), B1 => l074_n_81, B2 => y(2), ZN => l074_n_117);
  l074_g12552 : ND2D1BWP7T port map(A1 => l074_n_107, A2 => l074_n_2, ZN => l074_n_109);
  l074_g12553 : MAOI22D0BWP7T port map(A1 => l074_n_42, A2 => y(1), B1 => l074_n_42, B2 => y(1), ZN => l074_n_116);
  l074_g12554 : INR3D0BWP7T port map(A1 => l074_n_78, B1 => l074_n_62, B2 => l074_n_77, ZN => l074_n_115);
  l074_g12555 : MOAI22D0BWP7T port map(A1 => l074_n_47, A2 => y(0), B1 => l074_n_47, B2 => y(0), ZN => l074_n_114);
  l074_g12556 : MAOI22D0BWP7T port map(A1 => l074_n_41, A2 => l074_n_22, B1 => l074_n_41, B2 => l074_n_22, ZN => l074_n_113);
  l074_g12557 : MOAI22D0BWP7T port map(A1 => l074_n_41, A2 => l074_n_24, B1 => l074_n_41, B2 => l074_n_24, ZN => l074_n_112);
  l074_g12558 : NR2D0BWP7T port map(A1 => l074_n_46, A2 => l074_n_31, ZN => l074_n_100);
  l074_g12559 : NR2D1BWP7T port map(A1 => l074_n_46, A2 => l074_n_25, ZN => l074_n_99);
  l074_g12561 : AN2D1BWP7T port map(A1 => l074_n_52, A2 => l074_n_29, Z => l074_n_108);
  l074_g12562 : ND2D1BWP7T port map(A1 => l074_n_42, A2 => l074_n_32, ZN => l074_n_107);
  l074_g12563 : NR2D0BWP7T port map(A1 => l074_n_82, A2 => y_enemy4(5), ZN => l074_n_98);
  l074_g12564 : CKAN2D1BWP7T port map(A1 => l074_n_49, A2 => l074_n_39, Z => l074_n_106);
  l074_g12565 : ND2D1BWP7T port map(A1 => l074_n_67, A2 => l074_n_17, ZN => l074_n_105);
  l074_g12566 : OR2D1BWP7T port map(A1 => l074_n_49, A2 => l074_n_16, Z => l074_n_104);
  l074_g12567 : NR2XD0BWP7T port map(A1 => l074_n_67, A2 => l074_n_17, ZN => l074_n_97);
  l074_g12568 : CKAN2D1BWP7T port map(A1 => l074_n_15, A2 => l074_n_39, Z => l074_n_103);
  l074_g12569 : INR2D1BWP7T port map(A1 => l074_n_47, B1 => l074_n_45, ZN => l074_n_102);
  l074_g12570 : NR2XD0BWP7T port map(A1 => l074_n_72, A2 => l074_n_79, ZN => l074_n_101);
  l074_g12571 : NR2D0BWP7T port map(A1 => l074_n_53, A2 => l074_n_34, ZN => l074_n_89);
  l074_g12572 : AOI22D0BWP7T port map(A1 => l074_n_59, A2 => l074_n_13, B1 => l074_n_62, B2 => l074_n_26, ZN => l074_n_88);
  l074_g12573 : AOI22D0BWP7T port map(A1 => l074_n_54, A2 => x(0), B1 => x(1), B2 => l074_n_10, ZN => l074_n_87);
  l074_g12574 : AOI21D0BWP7T port map(A1 => l074_n_57, A2 => l074_n_60, B => draw_count8(1), ZN => l074_n_86);
  l074_g12575 : OA21D0BWP7T port map(A1 => l074_n_58, A2 => l074_n_55, B => l074_n_26, Z => l074_n_85);
  l074_g12576 : AOI21D0BWP7T port map(A1 => l074_n_58, A2 => l074_n_26, B => l074_n_63, ZN => l074_n_84);
  l074_g12577 : OAI21D0BWP7T port map(A1 => l074_n_56, A2 => draw_count8(1), B => l074_n_74, ZN => l074_n_96);
  l074_g12578 : AOI21D0BWP7T port map(A1 => l074_n_62, A2 => l074_n_12, B => l074_n_59, ZN => l074_n_95);
  l074_g12579 : OAI21D0BWP7T port map(A1 => l074_n_63, A2 => l074_n_55, B => l074_n_13, ZN => l074_n_94);
  l074_g12580 : MOAI22D0BWP7T port map(A1 => l074_n_0, A2 => l074_n_27, B1 => l074_n_66, B2 => l074_n_13, ZN => l074_n_93);
  l074_g12581 : AO21D0BWP7T port map(A1 => l074_n_64, A2 => l074_n_27, B => l074_n_72, Z => l074_n_92);
  l074_g12582 : IOA21D1BWP7T port map(A1 => l074_n_58, A2 => l074_n_12, B => l074_n_76, ZN => l074_n_91);
  l074_g12583 : OAI22D0BWP7T port map(A1 => l074_n_57, A2 => l074_n_12, B1 => l074_n_60, B2 => l074_n_27, ZN => l074_n_90);
  l074_g12584 : INVD1BWP7T port map(I => l074_n_42, ZN => l074_n_83);
  l074_g12586 : INVD1BWP7T port map(I => l074_n_48, ZN => l074_n_82);
  l074_g12587 : INVD0BWP7T port map(I => l074_n_41, ZN => l074_n_81);
  l074_g12588 : ND2D1BWP7T port map(A1 => l074_n_59, A2 => draw_count8(1), ZN => l074_n_80);
  l074_g12589 : NR2D1BWP7T port map(A1 => l074_n_0, A2 => draw_count8(1), ZN => l074_n_79);
  l074_g12590 : IND2D0BWP7T port map(A1 => l074_n_14, B1 => l074_n_63, ZN => l074_n_78);
  l074_g12591 : INR2D1BWP7T port map(A1 => l074_n_59, B1 => draw_count8(1), ZN => l074_n_77);
  l074_g12592 : CKND2D0BWP7T port map(A1 => l074_n_63, A2 => l074_n_13, ZN => l074_n_76);
  l074_g12593 : NR2D0BWP7T port map(A1 => l074_n_56, A2 => l074_n_7, ZN => l074_n_75);
  l074_g12594 : NR2D0BWP7T port map(A1 => l074_n_60, A2 => l074_n_14, ZN => l074_n_68);
  l074_g12595 : CKND2D1BWP7T port map(A1 => l074_n_58, A2 => l074_n_65, ZN => l074_n_74);
  l074_g12596 : IND2D1BWP7T port map(A1 => l074_n_59, B1 => l074_n_61, ZN => l074_n_73);
  l074_g12597 : AN2D0BWP7T port map(A1 => l074_n_63, A2 => l074_n_26, Z => l074_n_72);
  l074_g12598 : ND2D1BWP7T port map(A1 => l074_n_55, A2 => l074_n_12, ZN => l074_n_71);
  l074_g12599 : INR2D1BWP7T port map(A1 => l074_n_28, B1 => l074_n_57, ZN => l074_n_70);
  l074_g12600 : ND2D1BWP7T port map(A1 => l074_n_63, A2 => l074_n_65, ZN => l074_n_69);
  l074_g12601 : INVD1BWP7T port map(I => l074_n_0, ZN => l074_n_64);
  l074_g12602 : INVD1BWP7T port map(I => l074_n_62, ZN => l074_n_61);
  l074_g12603 : INVD0BWP7T port map(I => l074_n_58, ZN => l074_n_57);
  l074_g12604 : INVD1BWP7T port map(I => l074_n_56, ZN => l074_n_55);
  l074_g12605 : IAO21D0BWP7T port map(A1 => x(1), A2 => l074_n_10, B => x_enemy4(0), ZN => l074_n_54);
  l074_g12606 : AO21D0BWP7T port map(A1 => x(4), A2 => l074_n_11, B => l074_n_15, Z => l074_n_67);
  l074_g12607 : INR2D1BWP7T port map(A1 => draw_count8(3), B1 => l074_n_33, ZN => l074_n_66);
  l074_g12608 : IND2D1BWP7T port map(A1 => l074_n_28, B1 => l074_n_14, ZN => l074_n_65);
  l074_g12610 : NR2D1BWP7T port map(A1 => l074_n_33, A2 => draw_count8(3), ZN => l074_n_63);
  l074_g12611 : INR2D1BWP7T port map(A1 => l074_n_23, B1 => draw_count8(3), ZN => l074_n_62);
  l074_g12612 : ND2D1BWP7T port map(A1 => l074_n_37, A2 => draw_count8(3), ZN => l074_n_60);
  l074_g12613 : NR2D1BWP7T port map(A1 => l074_n_38, A2 => draw_count8(3), ZN => l074_n_59);
  l074_g12614 : NR2D1BWP7T port map(A1 => l074_n_40, A2 => draw_count8(3), ZN => l074_n_58);
  l074_g12615 : ND2D1BWP7T port map(A1 => l074_n_23, A2 => draw_count8(3), ZN => l074_n_56);
  l074_g12617 : INVD0BWP7T port map(I => l074_n_45, ZN => l074_n_44);
  l074_g12618 : MOAI22D0BWP7T port map(A1 => y(8), A2 => y_enemy4(8), B1 => y(8), B2 => y_enemy4(8), ZN => l074_n_53);
  l074_g12619 : MAOI22D0BWP7T port map(A1 => y(7), A2 => y_enemy4(7), B1 => y(7), B2 => y_enemy4(7), ZN => l074_n_52);
  l074_g12620 : MOAI22D0BWP7T port map(A1 => x(7), A2 => x_enemy4(7), B1 => x(7), B2 => x_enemy4(7), ZN => l074_n_51);
  l074_g12621 : MAOI22D0BWP7T port map(A1 => x(3), A2 => x_enemy4(3), B1 => x(3), B2 => x_enemy4(3), ZN => l074_n_50);
  l074_g12622 : MAOI22D0BWP7T port map(A1 => x(6), A2 => x_enemy4(6), B1 => x(6), B2 => x_enemy4(6), ZN => l074_n_49);
  l074_g12623 : OAI21D0BWP7T port map(A1 => l074_n_8, A2 => y_enemy4(6), B => l074_n_29, ZN => l074_n_48);
  l074_g12624 : MOAI22D0BWP7T port map(A1 => y(1), A2 => y_enemy4(1), B1 => y(1), B2 => y_enemy4(1), ZN => l074_n_47);
  l074_g12625 : MAOI22D0BWP7T port map(A1 => y(5), A2 => y_enemy4(5), B1 => y(5), B2 => y_enemy4(5), ZN => l074_n_46);
  l074_g12626 : MAOI22D0BWP7T port map(A1 => y(0), A2 => y_enemy4(0), B1 => y(0), B2 => y_enemy4(0), ZN => l074_n_45);
  l074_g12627 : MOAI22D0BWP7T port map(A1 => y(4), A2 => y_enemy4(4), B1 => y(4), B2 => y_enemy4(4), ZN => l074_n_43);
  l074_g12628 : MAOI22D0BWP7T port map(A1 => y(2), A2 => y_enemy4(2), B1 => y(2), B2 => y_enemy4(2), ZN => l074_n_42);
  l074_g12629 : MOAI22D0BWP7T port map(A1 => y(3), A2 => y_enemy4(3), B1 => y(3), B2 => y_enemy4(3), ZN => l074_n_41);
  l074_g12631 : CKND1BWP7T port map(I => l074_n_37, ZN => l074_n_38);
  l074_g12632 : INVD1BWP7T port map(I => l074_n_27, ZN => l074_n_26);
  l074_g12633 : IND2D1BWP7T port map(A1 => draw_count8(2), B1 => draw_count8(4), ZN => l074_n_40);
  l074_g12634 : IND2D1BWP7T port map(A1 => x_enemy4(5), B1 => x(5), ZN => l074_n_39);
  l074_g12635 : INR2D1BWP7T port map(A1 => draw_count8(2), B1 => draw_count8(4), ZN => l074_n_37);
  l074_g12636 : IND2D0BWP7T port map(A1 => y_enemy4(3), B1 => y(3), ZN => l074_n_36);
  l074_g12637 : IND2D0BWP7T port map(A1 => y_enemy4(1), B1 => y(1), ZN => l074_n_35);
  l074_g12638 : INR2XD0BWP7T port map(A1 => y_enemy4(7), B1 => y(7), ZN => l074_n_34);
  l074_g12639 : ND2D1BWP7T port map(A1 => draw_count8(2), A2 => draw_count8(4), ZN => l074_n_33);
  l074_g12640 : IND2D1BWP7T port map(A1 => y(1), B1 => y_enemy4(1), ZN => l074_n_32);
  l074_g12641 : IND2D1BWP7T port map(A1 => y_enemy4(4), B1 => y(4), ZN => l074_n_31);
  l074_g12642 : IND2D1BWP7T port map(A1 => x(7), B1 => x_enemy4(7), ZN => l074_n_30);
  l074_g12643 : ND2D1BWP7T port map(A1 => l074_n_8, A2 => y_enemy4(6), ZN => l074_n_29);
  l074_g12644 : INR2D1BWP7T port map(A1 => draw_count8(0), B1 => draw_count8(1), ZN => l074_n_28);
  l074_g12645 : CKND2D1BWP7T port map(A1 => draw_count8(1), A2 => draw_count8(0), ZN => l074_n_27);
  l074_g12646 : INVD1BWP7T port map(I => l074_n_13, ZN => l074_n_12);
  l074_g12647 : INR2XD0BWP7T port map(A1 => y_enemy4(4), B1 => y(4), ZN => l074_n_25);
  l074_g12648 : IND2D1BWP7T port map(A1 => y(2), B1 => y_enemy4(2), ZN => l074_n_24);
  l074_g12649 : NR2D0BWP7T port map(A1 => draw_count8(2), A2 => draw_count8(4), ZN => l074_n_23);
  l074_g12650 : IND2D1BWP7T port map(A1 => y_enemy4(2), B1 => y(2), ZN => l074_n_22);
  l074_g12651 : NR2D0BWP7T port map(A1 => l074_n_9, A2 => x_enemy4(8), ZN => l074_n_21);
  l074_g12652 : IND2D1BWP7T port map(A1 => y(8), B1 => y_enemy4(8), ZN => l074_n_20);
  l074_g12653 : IND2D1BWP7T port map(A1 => y(3), B1 => y_enemy4(3), ZN => l074_n_19);
  l074_g12654 : IND2D1BWP7T port map(A1 => x_enemy4(6), B1 => x(6), ZN => l074_n_18);
  l074_g12655 : IND2D1BWP7T port map(A1 => x(3), B1 => x_enemy4(3), ZN => l074_n_17);
  l074_g12656 : INR2XD0BWP7T port map(A1 => x_enemy4(5), B1 => x(5), ZN => l074_n_16);
  l074_g12657 : NR2D0BWP7T port map(A1 => x(4), A2 => l074_n_11, ZN => l074_n_15);
  l074_g12658 : IND2D1BWP7T port map(A1 => draw_count8(0), B1 => draw_count8(1), ZN => l074_n_14);
  l074_g12659 : NR2D0BWP7T port map(A1 => draw_count8(1), A2 => draw_count8(0), ZN => l074_n_13);
  l074_g12660 : CKND1BWP7T port map(I => x_enemy4(4), ZN => l074_n_11);
  l074_g12661 : INVD0BWP7T port map(I => x_enemy4(1), ZN => l074_n_10);
  l074_g12662 : CKND1BWP7T port map(I => x(8), ZN => l074_n_9);
  l074_g12663 : CKND1BWP7T port map(I => y(6), ZN => l074_n_8);
  l074_g12664 : INVD0BWP7T port map(I => draw_count8(1), ZN => l074_n_7);
  l074_g2 : INR3D0BWP7T port map(A1 => l074_n_121, B1 => l074_n_114, B2 => l074_n_44, ZN => l074_n_6);
  l074_g12665 : IND2D1BWP7T port map(A1 => l074_n_118, B1 => l074_n_175, ZN => l074_n_5);
  l074_g12666 : INR3D0BWP7T port map(A1 => l074_n_116, B1 => l074_n_45, B2 => l074_n_47, ZN => l074_n_4);
  l074_g12667 : IIND4D0BWP7T port map(A1 => l074_n_120, A2 => l074_n_112, B1 => l074_n_149, B2 => l074_n_176, ZN => l074_n_3);
  l074_g12668 : IND2D1BWP7T port map(A1 => l074_n_32, B1 => l074_n_83, ZN => l074_n_2);
  l074_g12669 : INR3D0BWP7T port map(A1 => l074_n_46, B1 => l074_n_133, B2 => l074_n_81, ZN => l074_n_1);
  l074_g12670 : IND2D1BWP7T port map(A1 => l074_n_40, B1 => draw_count8(3), ZN => l074_n_0);
  l03_hold_reg : DFD1BWP7T port map(CP => clk, D => l03_n_9, Q => UNCONNECTED, QN => l03_n_11);
  l03_g306 : INVD4BWP7T port map(I => l03_n_11, ZN => hsync);
  l03_g307 : INVD4BWP7T port map(I => l03_vold, ZN => vsync);
  l03_vold_reg : DFD1BWP7T port map(CP => clk, D => l03_n_0, Q => UNCONNECTED0, QN => l03_vold);
  l03_g309 : NR2XD0BWP7T port map(A1 => l03_n_33, A2 => reset, ZN => l03_n_9);
  l03_g312 : OAI21D0BWP7T port map(A1 => l03_n_4, A2 => x(8), B => l03_n_2, ZN => l03_n_7);
  l03_g313 : NR4D0BWP7T port map(A1 => l03_n_1, A2 => y(2), A3 => y(6), A4 => y(9), ZN => l03_n_6);
  l03_g314 : NR3D0BWP7T port map(A1 => x(6), A2 => x(4), A3 => x(5), ZN => l03_n_5);
  l03_g315 : AOI21D0BWP7T port map(A1 => x(4), A2 => x(5), B => x(6), ZN => l03_n_4);
  l03_g316 : NR4D0BWP7T port map(A1 => y(7), A2 => y(8), A3 => y(5), A4 => y(4), ZN => l03_n_3);
  l03_g317 : XNR2D1BWP7T port map(A1 => x(8), A2 => x(7), ZN => l03_n_2);
  l03_g318 : OR2D1BWP7T port map(A1 => y(1), A2 => y(3), Z => l03_n_1);
  l03_g2 : AOI21D0BWP7T port map(A1 => l03_n_6, A2 => l03_n_3, B => reset, ZN => l03_n_0);
  l03_g320 : AOI21D0BWP7T port map(A1 => l03_n_5, A2 => x(8), B => l03_n_7, ZN => l03_n_33);
  l075_g12411 : OAI221D0BWP7T port map(A1 => l075_n_221, A2 => l075_n_183, B1 => l075_n_155, B2 => l075_n_224, C => l075_n_245, ZN => r9);
  l075_g12412 : NR4D0BWP7T port map(A1 => l075_n_244, A2 => l075_n_234, A3 => l075_n_228, A4 => l075_n_205, ZN => l075_n_245);
  l075_g12413 : IND4D0BWP7T port map(A1 => l075_n_232, B1 => l075_n_227, B2 => l075_n_233, B3 => l075_n_241, ZN => l075_n_244);
  l075_g12414 : AO211D0BWP7T port map(A1 => l075_n_217, A2 => l075_n_91, B => l075_n_242, C => l075_n_240, Z => g9);
  l075_g12415 : OAI211D1BWP7T port map(A1 => l075_n_125, A2 => l075_n_221, B => l075_n_238, C => l075_n_230, ZN => l075_n_242);
  l075_g12416 : MAOI22D0BWP7T port map(A1 => l075_n_214, A2 => l075_n_161, B1 => l075_n_235, B2 => l075_n_193, ZN => l075_n_241);
  l075_g12417 : AO221D0BWP7T port map(A1 => l075_n_214, A2 => l075_n_138, B1 => l075_n_211, B2 => l075_n_126, C => l075_n_236, Z => l075_n_240);
  l075_g12418 : OAI32D0BWP7T port map(A1 => l075_n_26, A2 => l075_n_61, A3 => l075_n_221, B1 => l075_n_95, B2 => l075_n_223, ZN => b9);
  l075_g12419 : AOI211XD0BWP7T port map(A1 => l075_n_198, A2 => l075_n_70, B => l075_n_231, C => l075_n_225, ZN => l075_n_238);
  l075_g12420 : ND3D0BWP7T port map(A1 => l075_n_219, A2 => l075_n_210, A3 => l075_n_197, ZN => enable9);
  l075_g12421 : OAI211D1BWP7T port map(A1 => l075_n_84, A2 => l075_n_203, B => l075_n_218, C => l075_n_226, ZN => l075_n_236);
  l075_g12422 : ND4D0BWP7T port map(A1 => l075_n_215, A2 => l075_n_186, A3 => l075_n_180, A4 => l075_n_164, ZN => l075_n_235);
  l075_g12423 : OAI211D1BWP7T port map(A1 => l075_n_171, A2 => l075_n_223, B => l075_n_220, C => l075_n_206, ZN => l075_n_234);
  l075_g12424 : AOI22D0BWP7T port map(A1 => l075_n_211, A2 => l075_n_156, B1 => l075_n_216, B2 => l075_n_160, ZN => l075_n_233);
  l075_g12425 : AOI31D0BWP7T port map(A1 => l075_n_129, A2 => l075_n_131, A3 => l075_n_61, B => l075_n_229, ZN => l075_n_232);
  l075_g12426 : AOI21D0BWP7T port map(A1 => l075_n_131, A2 => l075_n_71, B => l075_n_224, ZN => l075_n_231);
  l075_g12427 : OAI21D0BWP7T port map(A1 => l075_n_132, A2 => l075_n_91, B => l075_n_222, ZN => l075_n_230);
  l075_g12428 : AOI21D0BWP7T port map(A1 => l075_n_209, A2 => l075_n_149, B => l075_n_195, ZN => l075_n_229);
  l075_g12429 : IAO21D0BWP7T port map(A1 => l075_n_152, A2 => l075_n_70, B => l075_n_212, ZN => l075_n_228);
  l075_g12430 : OAI31D0BWP7T port map(A1 => l075_n_75, A2 => l075_n_91, A3 => l075_n_111, B => l075_n_213, ZN => l075_n_227);
  l075_g12431 : OAI21D0BWP7T port map(A1 => l075_n_132, A2 => l075_n_138, B => l075_n_213, ZN => l075_n_226);
  l075_g12432 : AOI21D0BWP7T port map(A1 => l075_n_101, A2 => l075_n_69, B => l075_n_212, ZN => l075_n_225);
  l075_g12433 : CKND1BWP7T port map(I => l075_n_222, ZN => l075_n_223);
  l075_g12434 : OAI21D0BWP7T port map(A1 => l075_n_90, A2 => l075_n_55, B => l075_n_217, ZN => l075_n_220);
  l075_g12435 : AOI22D0BWP7T port map(A1 => l075_n_204, A2 => l075_n_192, B1 => l075_n_202, B2 => l075_n_177, ZN => l075_n_219);
  l075_g12436 : OAI21D0BWP7T port map(A1 => l075_n_92, A2 => l075_n_64, B => l075_n_216, ZN => l075_n_218);
  l075_g12437 : AOI22D0BWP7T port map(A1 => l075_n_208, A2 => l075_n_150, B1 => l075_n_209, B2 => l075_n_4, ZN => l075_n_224);
  l075_g12438 : OAI32D1BWP7T port map(A1 => l075_n_117, A2 => l075_n_134, A3 => l075_n_197, B1 => l075_n_157, B2 => l075_n_207, ZN => l075_n_222);
  l075_g12439 : AOI22D0BWP7T port map(A1 => l075_n_209, A2 => l075_n_6, B1 => l075_n_208, B2 => l075_n_151, ZN => l075_n_221);
  l075_g12440 : AOI211D1BWP7T port map(A1 => l075_n_127, A2 => l075_n_56, B => l075_n_196, C => l075_n_187, ZN => l075_n_215);
  l075_g12441 : OAI22D0BWP7T port map(A1 => l075_n_199, A2 => l075_n_170, B1 => l075_n_193, B2 => l075_n_180, ZN => l075_n_217);
  l075_g12442 : IOA21D1BWP7T port map(A1 => l075_n_202, A2 => l075_n_166, B => l075_n_210, ZN => l075_n_216);
  l075_g12443 : MOAI22D0BWP7T port map(A1 => l075_n_199, A2 => l075_n_164, B1 => l075_n_202, B2 => l075_n_165, ZN => l075_n_214);
  l075_g12444 : MOAI22D0BWP7T port map(A1 => l075_n_199, A2 => l075_n_167, B1 => l075_n_202, B2 => l075_n_168, ZN => l075_n_213);
  l075_g12445 : MAOI22D0BWP7T port map(A1 => l075_n_200, A2 => l075_n_165, B1 => l075_n_201, B2 => l075_n_164, ZN => l075_n_212);
  l075_g12446 : MOAI22D0BWP7T port map(A1 => l075_n_193, A2 => l075_n_186, B1 => l075_n_200, B2 => l075_n_166, ZN => l075_n_211);
  l075_g12447 : INVD0BWP7T port map(I => l075_n_208, ZN => l075_n_207);
  l075_g12448 : ND2D1BWP7T port map(A1 => l075_n_200, A2 => l075_n_148, ZN => l075_n_210);
  l075_g12449 : NR2D1BWP7T port map(A1 => l075_n_197, A2 => l075_n_112, ZN => l075_n_209);
  l075_g12450 : NR2D1BWP7T port map(A1 => l075_n_197, A2 => l075_n_113, ZN => l075_n_208);
  l075_g12451 : OAI21D0BWP7T port map(A1 => l075_n_130, A2 => l075_n_75, B => l075_n_198, ZN => l075_n_206);
  l075_g12452 : AOI21D0BWP7T port map(A1 => l075_n_142, A2 => l075_n_80, B => l075_n_203, ZN => l075_n_205);
  l075_g12453 : ND4D0BWP7T port map(A1 => l075_n_194, A2 => l075_n_189, A3 => l075_n_3, A4 => l075_n_181, ZN => l075_n_204);
  l075_g12454 : INVD0BWP7T port map(I => l075_n_202, ZN => l075_n_201);
  l075_g12455 : INVD0BWP7T port map(I => l075_n_200, ZN => l075_n_199);
  l075_g12456 : CKND2D1BWP7T port map(A1 => l075_n_192, A2 => l075_n_187, ZN => l075_n_203);
  l075_g12457 : NR2D1BWP7T port map(A1 => l075_n_193, A2 => l075_n_5, ZN => l075_n_202);
  l075_g12458 : NR2D1BWP7T port map(A1 => l075_n_193, A2 => l075_n_184, ZN => l075_n_200);
  l075_g12459 : OA31D1BWP7T port map(A1 => l075_n_119, A2 => l075_n_147, A3 => l075_n_174, B => l075_n_194, Z => l075_n_196);
  l075_g12460 : NR4D0BWP7T port map(A1 => l075_n_193, A2 => l075_n_172, A3 => l075_n_163, A4 => l075_n_43, ZN => l075_n_195);
  l075_g12461 : AOI21D0BWP7T port map(A1 => l075_n_3, A2 => l075_n_181, B => l075_n_193, ZN => l075_n_198);
  l075_g12462 : ND3D0BWP7T port map(A1 => l075_n_192, A2 => l075_n_175, A3 => l075_n_120, ZN => l075_n_197);
  l075_g12463 : INR2XD0BWP7T port map(A1 => l075_n_186, B1 => l075_n_191, ZN => l075_n_194);
  l075_g12464 : INVD1BWP7T port map(I => l075_n_193, ZN => l075_n_192);
  l075_g12465 : OAI221D0BWP7T port map(A1 => l075_n_173, A2 => l075_n_141, B1 => l075_n_30, B2 => l075_n_21, C => l075_n_190, ZN => l075_n_193);
  l075_g12466 : OAI221D0BWP7T port map(A1 => l075_n_184, A2 => l075_n_178, B1 => l075_n_170, B2 => l075_n_5, C => l075_n_180, ZN => l075_n_191);
  l075_g12467 : AOI221D0BWP7T port map(A1 => l075_n_9, A2 => x_enemy5(8), B1 => l075_n_51, B2 => l075_n_18, C => l075_n_185, ZN => l075_n_190);
  l075_g12468 : IAO21D0BWP7T port map(A1 => l075_n_5, A2 => l075_n_182, B => l075_n_188, ZN => l075_n_189);
  l075_g12469 : AOI21D0BWP7T port map(A1 => l075_n_182, A2 => l075_n_170, B => l075_n_184, ZN => l075_n_188);
  l075_g12470 : OAI22D0BWP7T port map(A1 => l075_n_5, A2 => l075_n_167, B1 => l075_n_184, B2 => l075_n_169, ZN => l075_n_187);
  l075_g12471 : IND2D1BWP7T port map(A1 => l075_n_5, B1 => l075_n_148, ZN => l075_n_186);
  l075_g12472 : AO21D0BWP7T port map(A1 => l075_n_21, A2 => l075_n_30, B => l075_n_179, Z => l075_n_185);
  l075_g12474 : NR3D0BWP7T port map(A1 => l075_n_162, A2 => l075_n_90, A3 => l075_n_64, ZN => l075_n_183);
  l075_g12475 : ND2D1BWP7T port map(A1 => l075_n_175, A2 => l075_n_118, ZN => l075_n_184);
  l075_g12477 : MOAI22D0BWP7T port map(A1 => l075_n_51, A2 => l075_n_18, B1 => l075_n_159, B2 => l075_n_141, ZN => l075_n_179);
  l075_g12478 : INR3D0BWP7T port map(A1 => l075_n_167, B1 => l075_n_165, B2 => l075_n_166, ZN => l075_n_182);
  l075_g12479 : ND4D0BWP7T port map(A1 => l075_n_1, A2 => l075_n_154, A3 => l075_n_145, A4 => l075_n_43, ZN => l075_n_181);
  l075_g12480 : IND3D1BWP7T port map(A1 => l075_n_147, B1 => l075_n_119, B2 => l075_n_176, ZN => l075_n_180);
  l075_g12481 : CKND1BWP7T port map(I => l075_n_177, ZN => l075_n_178);
  l075_g12482 : INVD0BWP7T port map(I => l075_n_175, ZN => l075_n_174);
  l075_g12483 : ND2D1BWP7T port map(A1 => l075_n_169, A2 => l075_n_164, ZN => l075_n_177);
  l075_g12484 : AOI211XD0BWP7T port map(A1 => l075_n_46, A2 => l075_n_31, B => l075_n_163, C => l075_n_100, ZN => l075_n_176);
  l075_g12485 : AOI211XD0BWP7T port map(A1 => l075_n_46, A2 => l075_n_25, B => l075_n_163, C => l075_n_99, ZN => l075_n_175);
  l075_g12486 : AOI221D0BWP7T port map(A1 => l075_n_106, A2 => l075_n_16, B1 => l075_n_49, B2 => l075_n_103, C => l075_n_158, ZN => l075_n_173);
  l075_g12487 : AOI22D0BWP7T port map(A1 => l075_n_1, A2 => y(4), B1 => l075_n_153, B2 => l075_n_41, ZN => l075_n_172);
  l075_g12488 : INR4D0BWP7T port map(A1 => l075_n_95, B1 => l075_n_93, B2 => l075_n_146, B3 => l075_n_132, ZN => l075_n_171);
  l075_g12489 : INVD0BWP7T port map(I => l075_n_169, ZN => l075_n_168);
  l075_g12490 : ND2D1BWP7T port map(A1 => l075_n_149, A2 => l075_n_112, ZN => l075_n_170);
  l075_g12491 : ND2D1BWP7T port map(A1 => l075_n_4, A2 => l075_n_112, ZN => l075_n_169);
  l075_g12492 : ND2D1BWP7T port map(A1 => l075_n_150, A2 => l075_n_113, ZN => l075_n_167);
  l075_g12493 : INR2D1BWP7T port map(A1 => l075_n_113, B1 => l075_n_157, ZN => l075_n_166);
  l075_g12494 : AN2D1BWP7T port map(A1 => l075_n_6, A2 => l075_n_112, Z => l075_n_165);
  l075_g12495 : ND2D1BWP7T port map(A1 => l075_n_151, A2 => l075_n_113, ZN => l075_n_164);
  l075_g12496 : IND4D0BWP7T port map(A1 => l075_n_70, B1 => l075_n_71, B2 => l075_n_101, B3 => l075_n_115, ZN => l075_n_162);
  l075_g12497 : ND4D0BWP7T port map(A1 => l075_n_128, A2 => l075_n_94, A3 => l075_n_69, A4 => l075_n_60, ZN => l075_n_161);
  l075_g12498 : IND4D0BWP7T port map(A1 => l075_n_75, B1 => l075_n_69, B2 => l075_n_76, B3 => l075_n_123, ZN => l075_n_160);
  l075_g12499 : OAI222D0BWP7T port map(A1 => l075_n_144, A2 => l075_n_137, B1 => l075_n_97, B2 => l075_n_136, C1 => l075_n_103, C2 => l075_n_104, ZN => l075_n_159);
  l075_g12500 : MOAI22D0BWP7T port map(A1 => l075_n_143, A2 => l075_n_135, B1 => l075_n_137, B2 => l075_n_105, ZN => l075_n_158);
  l075_g12501 : ND3D0BWP7T port map(A1 => l075_n_139, A2 => l075_n_145, A3 => l075_n_140, ZN => l075_n_163);
  l075_g12502 : OAI211D1BWP7T port map(A1 => l075_n_14, A2 => l075_n_56, B => l075_n_142, C => l075_n_88, ZN => l075_n_156);
  l075_g12503 : INR3D0BWP7T port map(A1 => l075_n_115, B1 => l075_n_92, B2 => l075_n_124, ZN => l075_n_155);
  l075_g12504 : AOI211D1BWP7T port map(A1 => l075_n_48, A2 => y(5), B => l075_n_122, C => l075_n_107, ZN => l075_n_154);
  l075_g12505 : NR3D0BWP7T port map(A1 => l075_n_133, A2 => l075_n_46, A3 => y(4), ZN => l075_n_153);
  l075_g12506 : AO211D0BWP7T port map(A1 => l075_n_59, A2 => l075_n_12, B => l075_n_146, C => l075_n_85, Z => l075_n_152);
  l075_g12507 : ND3D0BWP7T port map(A1 => l075_n_114, A2 => l075_n_109, A3 => l075_n_45, ZN => l075_n_157);
  l075_g12510 : NR3D0BWP7T port map(A1 => l075_n_116, A2 => l075_n_45, A3 => l075_n_47, ZN => l075_n_151);
  l075_g12512 : NR3D0BWP7T port map(A1 => l075_n_121, A2 => l075_n_114, A3 => l075_n_44, ZN => l075_n_150);
  l075_g12513 : AN4D1BWP7T port map(A1 => l075_n_114, A2 => l075_n_2, A3 => l075_n_108, A4 => l075_n_45, Z => l075_n_149);
  l075_g12514 : INR2D1BWP7T port map(A1 => l075_n_117, B1 => l075_n_134, ZN => l075_n_148);
  l075_g12515 : OR2D1BWP7T port map(A1 => l075_n_133, A2 => l075_n_41, Z => l075_n_147);
  l075_g12516 : ND2D1BWP7T port map(A1 => l075_n_131, A2 => l075_n_94, ZN => l075_n_146);
  l075_g12517 : AOI211XD0BWP7T port map(A1 => l075_n_53, A2 => l075_n_34, B => l075_n_89, C => l075_n_110, ZN => l075_n_145);
  l075_g12518 : CKND1BWP7T port map(I => l075_n_143, ZN => l075_n_144);
  l075_g12519 : AOI22D0BWP7T port map(A1 => l075_n_98, A2 => y(5), B1 => l075_n_82, B2 => y_enemy5(5), ZN => l075_n_140);
  l075_g12520 : NR2XD0BWP7T port map(A1 => l075_n_122, A2 => l075_n_107, ZN => l075_n_139);
  l075_g12521 : MAOI222D1BWP7T port map(A => l075_n_87, B => x(2), C => x_enemy5(2), ZN => l075_n_143);
  l075_g12522 : NR3D0BWP7T port map(A1 => l075_n_96, A2 => l075_n_90, A3 => l075_n_68, ZN => l075_n_142);
  l075_g12523 : OAI21D0BWP7T port map(A1 => l075_n_106, A2 => l075_n_15, B => l075_n_104, ZN => l075_n_141);
  l075_g12524 : CKND1BWP7T port map(I => l075_n_135, ZN => l075_n_136);
  l075_g12525 : INVD0BWP7T port map(I => l075_n_131, ZN => l075_n_130);
  l075_g12526 : AOI211XD0BWP7T port map(A1 => l075_n_59, A2 => l075_n_26, B => l075_n_96, C => l075_n_79, ZN => l075_n_129);
  l075_g12527 : OAI21D0BWP7T port map(A1 => l075_n_73, A2 => l075_n_58, B => draw_count9(1), ZN => l075_n_128);
  l075_g12528 : AOI221D0BWP7T port map(A1 => l075_n_58, A2 => l075_n_27, B1 => l075_n_62, B2 => draw_count9(0), C => l075_n_77, ZN => l075_n_127);
  l075_g12529 : AO221D0BWP7T port map(A1 => l075_n_65, A2 => l075_n_64, B1 => l075_n_66, B2 => l075_n_28, C => l075_n_93, Z => l075_n_126);
  l075_g12530 : OA211D0BWP7T port map(A1 => l075_n_26, A2 => l075_n_60, B => l075_n_101, C => l075_n_78, Z => l075_n_125);
  l075_g12531 : OAI211D1BWP7T port map(A1 => l075_n_12, A2 => l075_n_56, B => l075_n_80, C => l075_n_74, ZN => l075_n_124);
  l075_g12532 : AOI21D0BWP7T port map(A1 => l075_n_59, A2 => l075_n_27, B => l075_n_86, ZN => l075_n_123);
  l075_g12533 : AO21D0BWP7T port map(A1 => l075_n_66, A2 => l075_n_65, B => l075_n_93, Z => l075_n_138);
  l075_g12534 : OAI22D0BWP7T port map(A1 => l075_n_67, A2 => l075_n_17, B1 => l075_n_50, B2 => x(2), ZN => l075_n_137);
  l075_g12535 : IOA21D1BWP7T port map(A1 => l075_n_50, A2 => x(2), B => l075_n_105, ZN => l075_n_135);
  l075_g12536 : ND2D1BWP7T port map(A1 => l075_n_102, A2 => l075_n_42, ZN => l075_n_134);
  l075_g12537 : ND2D1BWP7T port map(A1 => l075_n_102, A2 => l075_n_83, ZN => l075_n_133);
  l075_g12538 : IND2D1BWP7T port map(A1 => l075_n_92, B1 => l075_n_69, ZN => l075_n_132);
  l075_g12539 : INR2XD0BWP7T port map(A1 => l075_n_60, B1 => l075_n_90, ZN => l075_n_131);
  l075_g12544 : OAI22D0BWP7T port map(A1 => l075_n_52, A2 => l075_n_29, B1 => l075_n_48, B2 => y(5), ZN => l075_n_122);
  l075_g12545 : MOAI22D0BWP7T port map(A1 => l075_n_60, A2 => draw_count9(1), B1 => l075_n_73, B2 => l075_n_65, ZN => l075_n_111);
  l075_g12546 : MOAI22D0BWP7T port map(A1 => l075_n_20, A2 => y(9), B1 => l075_n_20, B2 => y(9), ZN => l075_n_110);
  l075_g12547 : MAOI22D0BWP7T port map(A1 => l075_n_83, A2 => l075_n_35, B1 => l075_n_83, B2 => l075_n_35, ZN => l075_n_121);
  l075_g12548 : MAOI22D0BWP7T port map(A1 => l075_n_43, A2 => l075_n_36, B1 => l075_n_43, B2 => l075_n_36, ZN => l075_n_120);
  l075_g12549 : MAOI22D0BWP7T port map(A1 => l075_n_43, A2 => y(3), B1 => l075_n_43, B2 => y(3), ZN => l075_n_119);
  l075_g12550 : MOAI22D0BWP7T port map(A1 => l075_n_43, A2 => l075_n_19, B1 => l075_n_43, B2 => l075_n_19, ZN => l075_n_118);
  l075_g12551 : MAOI22D0BWP7T port map(A1 => l075_n_81, A2 => y(2), B1 => l075_n_81, B2 => y(2), ZN => l075_n_117);
  l075_g12552 : ND2D1BWP7T port map(A1 => l075_n_2, A2 => l075_n_108, ZN => l075_n_109);
  l075_g12553 : MAOI22D0BWP7T port map(A1 => l075_n_42, A2 => y(1), B1 => l075_n_42, B2 => y(1), ZN => l075_n_116);
  l075_g12554 : INR3D0BWP7T port map(A1 => l075_n_78, B1 => l075_n_62, B2 => l075_n_77, ZN => l075_n_115);
  l075_g12555 : MOAI22D0BWP7T port map(A1 => l075_n_47, A2 => y(0), B1 => l075_n_47, B2 => y(0), ZN => l075_n_114);
  l075_g12556 : MAOI22D0BWP7T port map(A1 => l075_n_41, A2 => l075_n_22, B1 => l075_n_41, B2 => l075_n_22, ZN => l075_n_113);
  l075_g12557 : MOAI22D0BWP7T port map(A1 => l075_n_41, A2 => l075_n_24, B1 => l075_n_41, B2 => l075_n_24, ZN => l075_n_112);
  l075_g12558 : NR2XD0BWP7T port map(A1 => l075_n_46, A2 => l075_n_31, ZN => l075_n_100);
  l075_g12559 : NR2XD0BWP7T port map(A1 => l075_n_46, A2 => l075_n_25, ZN => l075_n_99);
  l075_g12560 : ND2D1BWP7T port map(A1 => l075_n_83, A2 => l075_n_32, ZN => l075_n_108);
  l075_g12561 : AN2D1BWP7T port map(A1 => l075_n_52, A2 => l075_n_29, Z => l075_n_107);
  l075_g12563 : NR2D0BWP7T port map(A1 => l075_n_82, A2 => y_enemy5(5), ZN => l075_n_98);
  l075_g12564 : CKAN2D1BWP7T port map(A1 => l075_n_49, A2 => l075_n_39, Z => l075_n_106);
  l075_g12565 : ND2D1BWP7T port map(A1 => l075_n_67, A2 => l075_n_17, ZN => l075_n_105);
  l075_g12566 : OR2D1BWP7T port map(A1 => l075_n_49, A2 => l075_n_16, Z => l075_n_104);
  l075_g12567 : NR2XD0BWP7T port map(A1 => l075_n_67, A2 => l075_n_17, ZN => l075_n_97);
  l075_g12568 : CKAN2D1BWP7T port map(A1 => l075_n_15, A2 => l075_n_39, Z => l075_n_103);
  l075_g12569 : INR2D1BWP7T port map(A1 => l075_n_47, B1 => l075_n_45, ZN => l075_n_102);
  l075_g12570 : NR2XD0BWP7T port map(A1 => l075_n_72, A2 => l075_n_79, ZN => l075_n_101);
  l075_g12571 : NR2D0BWP7T port map(A1 => l075_n_53, A2 => l075_n_34, ZN => l075_n_89);
  l075_g12572 : AOI22D0BWP7T port map(A1 => l075_n_59, A2 => l075_n_13, B1 => l075_n_62, B2 => l075_n_26, ZN => l075_n_88);
  l075_g12573 : AOI22D0BWP7T port map(A1 => l075_n_54, A2 => x(0), B1 => x(1), B2 => l075_n_10, ZN => l075_n_87);
  l075_g12574 : AOI21D0BWP7T port map(A1 => l075_n_57, A2 => l075_n_60, B => draw_count9(1), ZN => l075_n_86);
  l075_g12575 : OA21D0BWP7T port map(A1 => l075_n_58, A2 => l075_n_55, B => l075_n_26, Z => l075_n_85);
  l075_g12576 : AOI21D0BWP7T port map(A1 => l075_n_58, A2 => l075_n_26, B => l075_n_63, ZN => l075_n_84);
  l075_g12577 : OAI21D0BWP7T port map(A1 => l075_n_56, A2 => draw_count9(1), B => l075_n_74, ZN => l075_n_96);
  l075_g12578 : AOI21D0BWP7T port map(A1 => l075_n_62, A2 => l075_n_12, B => l075_n_59, ZN => l075_n_95);
  l075_g12579 : OAI21D0BWP7T port map(A1 => l075_n_63, A2 => l075_n_55, B => l075_n_13, ZN => l075_n_94);
  l075_g12580 : MOAI22D0BWP7T port map(A1 => l075_n_0, A2 => l075_n_27, B1 => l075_n_66, B2 => l075_n_13, ZN => l075_n_93);
  l075_g12581 : AO21D0BWP7T port map(A1 => l075_n_64, A2 => l075_n_27, B => l075_n_72, Z => l075_n_92);
  l075_g12582 : IOA21D1BWP7T port map(A1 => l075_n_58, A2 => l075_n_12, B => l075_n_76, ZN => l075_n_91);
  l075_g12583 : OAI22D0BWP7T port map(A1 => l075_n_57, A2 => l075_n_12, B1 => l075_n_60, B2 => l075_n_27, ZN => l075_n_90);
  l075_g12584 : INVD1BWP7T port map(I => l075_n_42, ZN => l075_n_83);
  l075_g12586 : INVD0BWP7T port map(I => l075_n_48, ZN => l075_n_82);
  l075_g12587 : INVD0BWP7T port map(I => l075_n_41, ZN => l075_n_81);
  l075_g12588 : ND2D1BWP7T port map(A1 => l075_n_59, A2 => draw_count9(1), ZN => l075_n_80);
  l075_g12589 : NR2D1BWP7T port map(A1 => l075_n_0, A2 => draw_count9(1), ZN => l075_n_79);
  l075_g12590 : IND2D0BWP7T port map(A1 => l075_n_14, B1 => l075_n_63, ZN => l075_n_78);
  l075_g12591 : INR2D1BWP7T port map(A1 => l075_n_59, B1 => draw_count9(1), ZN => l075_n_77);
  l075_g12592 : CKND2D0BWP7T port map(A1 => l075_n_63, A2 => l075_n_13, ZN => l075_n_76);
  l075_g12593 : NR2D0BWP7T port map(A1 => l075_n_56, A2 => l075_n_7, ZN => l075_n_75);
  l075_g12594 : NR2D0BWP7T port map(A1 => l075_n_60, A2 => l075_n_14, ZN => l075_n_68);
  l075_g12595 : CKND2D1BWP7T port map(A1 => l075_n_58, A2 => l075_n_65, ZN => l075_n_74);
  l075_g12596 : IND2D1BWP7T port map(A1 => l075_n_59, B1 => l075_n_61, ZN => l075_n_73);
  l075_g12597 : AN2D0BWP7T port map(A1 => l075_n_63, A2 => l075_n_26, Z => l075_n_72);
  l075_g12598 : ND2D1BWP7T port map(A1 => l075_n_55, A2 => l075_n_12, ZN => l075_n_71);
  l075_g12599 : INR2D1BWP7T port map(A1 => l075_n_28, B1 => l075_n_57, ZN => l075_n_70);
  l075_g12600 : ND2D1BWP7T port map(A1 => l075_n_63, A2 => l075_n_65, ZN => l075_n_69);
  l075_g12601 : INVD1BWP7T port map(I => l075_n_0, ZN => l075_n_64);
  l075_g12602 : INVD0BWP7T port map(I => l075_n_62, ZN => l075_n_61);
  l075_g12603 : INVD0BWP7T port map(I => l075_n_58, ZN => l075_n_57);
  l075_g12604 : INVD1BWP7T port map(I => l075_n_56, ZN => l075_n_55);
  l075_g12605 : IAO21D0BWP7T port map(A1 => x(1), A2 => l075_n_10, B => x_enemy5(0), ZN => l075_n_54);
  l075_g12606 : AO21D0BWP7T port map(A1 => x(4), A2 => l075_n_11, B => l075_n_15, Z => l075_n_67);
  l075_g12607 : INR2D1BWP7T port map(A1 => draw_count9(3), B1 => l075_n_33, ZN => l075_n_66);
  l075_g12608 : IND2D1BWP7T port map(A1 => l075_n_28, B1 => l075_n_14, ZN => l075_n_65);
  l075_g12610 : NR2D1BWP7T port map(A1 => l075_n_33, A2 => draw_count9(3), ZN => l075_n_63);
  l075_g12611 : INR2D1BWP7T port map(A1 => l075_n_23, B1 => draw_count9(3), ZN => l075_n_62);
  l075_g12612 : ND2D1BWP7T port map(A1 => l075_n_37, A2 => draw_count9(3), ZN => l075_n_60);
  l075_g12613 : NR2D1BWP7T port map(A1 => l075_n_38, A2 => draw_count9(3), ZN => l075_n_59);
  l075_g12614 : NR2D1BWP7T port map(A1 => l075_n_40, A2 => draw_count9(3), ZN => l075_n_58);
  l075_g12615 : ND2D1BWP7T port map(A1 => l075_n_23, A2 => draw_count9(3), ZN => l075_n_56);
  l075_g12617 : INVD0BWP7T port map(I => l075_n_45, ZN => l075_n_44);
  l075_g12618 : MOAI22D0BWP7T port map(A1 => y(8), A2 => y_enemy5(8), B1 => y(8), B2 => y_enemy5(8), ZN => l075_n_53);
  l075_g12619 : MAOI22D0BWP7T port map(A1 => y(7), A2 => y_enemy5(7), B1 => y(7), B2 => y_enemy5(7), ZN => l075_n_52);
  l075_g12620 : MOAI22D0BWP7T port map(A1 => x(7), A2 => x_enemy5(7), B1 => x(7), B2 => x_enemy5(7), ZN => l075_n_51);
  l075_g12621 : MAOI22D0BWP7T port map(A1 => x(3), A2 => x_enemy5(3), B1 => x(3), B2 => x_enemy5(3), ZN => l075_n_50);
  l075_g12622 : MAOI22D0BWP7T port map(A1 => x(6), A2 => x_enemy5(6), B1 => x(6), B2 => x_enemy5(6), ZN => l075_n_49);
  l075_g12623 : OAI21D0BWP7T port map(A1 => l075_n_8, A2 => y_enemy5(6), B => l075_n_29, ZN => l075_n_48);
  l075_g12624 : MOAI22D0BWP7T port map(A1 => y(1), A2 => y_enemy5(1), B1 => y(1), B2 => y_enemy5(1), ZN => l075_n_47);
  l075_g12625 : MAOI22D0BWP7T port map(A1 => y(5), A2 => y_enemy5(5), B1 => y(5), B2 => y_enemy5(5), ZN => l075_n_46);
  l075_g12626 : MAOI22D0BWP7T port map(A1 => y(0), A2 => y_enemy5(0), B1 => y(0), B2 => y_enemy5(0), ZN => l075_n_45);
  l075_g12627 : MOAI22D0BWP7T port map(A1 => y(4), A2 => y_enemy5(4), B1 => y(4), B2 => y_enemy5(4), ZN => l075_n_43);
  l075_g12628 : MAOI22D0BWP7T port map(A1 => y(2), A2 => y_enemy5(2), B1 => y(2), B2 => y_enemy5(2), ZN => l075_n_42);
  l075_g12629 : MOAI22D0BWP7T port map(A1 => y(3), A2 => y_enemy5(3), B1 => y(3), B2 => y_enemy5(3), ZN => l075_n_41);
  l075_g12631 : CKND1BWP7T port map(I => l075_n_37, ZN => l075_n_38);
  l075_g12632 : INVD1BWP7T port map(I => l075_n_27, ZN => l075_n_26);
  l075_g12633 : IND2D1BWP7T port map(A1 => draw_count9(2), B1 => draw_count9(4), ZN => l075_n_40);
  l075_g12634 : IND2D1BWP7T port map(A1 => x_enemy5(5), B1 => x(5), ZN => l075_n_39);
  l075_g12635 : INR2D1BWP7T port map(A1 => draw_count9(2), B1 => draw_count9(4), ZN => l075_n_37);
  l075_g12636 : IND2D0BWP7T port map(A1 => y_enemy5(3), B1 => y(3), ZN => l075_n_36);
  l075_g12637 : IND2D1BWP7T port map(A1 => y_enemy5(1), B1 => y(1), ZN => l075_n_35);
  l075_g12638 : INR2XD0BWP7T port map(A1 => y_enemy5(7), B1 => y(7), ZN => l075_n_34);
  l075_g12639 : ND2D1BWP7T port map(A1 => draw_count9(2), A2 => draw_count9(4), ZN => l075_n_33);
  l075_g12640 : INR2XD0BWP7T port map(A1 => y_enemy5(1), B1 => y(1), ZN => l075_n_32);
  l075_g12641 : IND2D1BWP7T port map(A1 => y_enemy5(4), B1 => y(4), ZN => l075_n_31);
  l075_g12642 : IND2D1BWP7T port map(A1 => x(7), B1 => x_enemy5(7), ZN => l075_n_30);
  l075_g12643 : ND2D1BWP7T port map(A1 => l075_n_8, A2 => y_enemy5(6), ZN => l075_n_29);
  l075_g12644 : INR2D1BWP7T port map(A1 => draw_count9(0), B1 => draw_count9(1), ZN => l075_n_28);
  l075_g12645 : CKND2D1BWP7T port map(A1 => draw_count9(1), A2 => draw_count9(0), ZN => l075_n_27);
  l075_g12646 : INVD1BWP7T port map(I => l075_n_13, ZN => l075_n_12);
  l075_g12647 : INR2XD0BWP7T port map(A1 => y_enemy5(4), B1 => y(4), ZN => l075_n_25);
  l075_g12648 : IND2D1BWP7T port map(A1 => y(2), B1 => y_enemy5(2), ZN => l075_n_24);
  l075_g12649 : NR2D0BWP7T port map(A1 => draw_count9(2), A2 => draw_count9(4), ZN => l075_n_23);
  l075_g12650 : IND2D1BWP7T port map(A1 => y_enemy5(2), B1 => y(2), ZN => l075_n_22);
  l075_g12651 : NR2D0BWP7T port map(A1 => l075_n_9, A2 => x_enemy5(8), ZN => l075_n_21);
  l075_g12652 : IND2D1BWP7T port map(A1 => y(8), B1 => y_enemy5(8), ZN => l075_n_20);
  l075_g12653 : IND2D1BWP7T port map(A1 => y(3), B1 => y_enemy5(3), ZN => l075_n_19);
  l075_g12654 : IND2D1BWP7T port map(A1 => x_enemy5(6), B1 => x(6), ZN => l075_n_18);
  l075_g12655 : IND2D1BWP7T port map(A1 => x(3), B1 => x_enemy5(3), ZN => l075_n_17);
  l075_g12656 : INR2XD0BWP7T port map(A1 => x_enemy5(5), B1 => x(5), ZN => l075_n_16);
  l075_g12657 : NR2D0BWP7T port map(A1 => x(4), A2 => l075_n_11, ZN => l075_n_15);
  l075_g12658 : IND2D1BWP7T port map(A1 => draw_count9(0), B1 => draw_count9(1), ZN => l075_n_14);
  l075_g12659 : NR2D0BWP7T port map(A1 => draw_count9(1), A2 => draw_count9(0), ZN => l075_n_13);
  l075_g12660 : CKND1BWP7T port map(I => x_enemy5(4), ZN => l075_n_11);
  l075_g12661 : INVD0BWP7T port map(I => x_enemy5(1), ZN => l075_n_10);
  l075_g12662 : CKND1BWP7T port map(I => x(8), ZN => l075_n_9);
  l075_g12663 : CKND1BWP7T port map(I => y(6), ZN => l075_n_8);
  l075_g12664 : INVD0BWP7T port map(I => draw_count9(1), ZN => l075_n_7);
  l075_g2 : INR3D0BWP7T port map(A1 => l075_n_121, B1 => l075_n_114, B2 => l075_n_44, ZN => l075_n_6);
  l075_g12665 : IND2D1BWP7T port map(A1 => l075_n_118, B1 => l075_n_176, ZN => l075_n_5);
  l075_g12666 : INR3D0BWP7T port map(A1 => l075_n_116, B1 => l075_n_45, B2 => l075_n_47, ZN => l075_n_4);
  l075_g12667 : IIND4D0BWP7T port map(A1 => l075_n_120, A2 => l075_n_112, B1 => l075_n_149, B2 => l075_n_176, ZN => l075_n_3);
  l075_g12668 : IND2D1BWP7T port map(A1 => l075_n_32, B1 => l075_n_42, ZN => l075_n_2);
  l075_g12669 : INR3D0BWP7T port map(A1 => l075_n_46, B1 => l075_n_133, B2 => l075_n_81, ZN => l075_n_1);
  l075_g12670 : IND2D1BWP7T port map(A1 => l075_n_40, B1 => draw_count9(3), ZN => l075_n_0);
  l076_g12411 : OAI221D0BWP7T port map(A1 => l076_n_221, A2 => l076_n_183, B1 => l076_n_155, B2 => l076_n_224, C => l076_n_245, ZN => r10);
  l076_g12412 : NR4D0BWP7T port map(A1 => l076_n_244, A2 => l076_n_234, A3 => l076_n_228, A4 => l076_n_205, ZN => l076_n_245);
  l076_g12413 : IND4D0BWP7T port map(A1 => l076_n_232, B1 => l076_n_227, B2 => l076_n_233, B3 => l076_n_241, ZN => l076_n_244);
  l076_g12414 : AO211D0BWP7T port map(A1 => l076_n_217, A2 => l076_n_91, B => l076_n_242, C => l076_n_240, Z => g10);
  l076_g12415 : OAI211D1BWP7T port map(A1 => l076_n_125, A2 => l076_n_221, B => l076_n_238, C => l076_n_230, ZN => l076_n_242);
  l076_g12416 : MAOI22D0BWP7T port map(A1 => l076_n_214, A2 => l076_n_161, B1 => l076_n_235, B2 => l076_n_193, ZN => l076_n_241);
  l076_g12417 : AO221D0BWP7T port map(A1 => l076_n_214, A2 => l076_n_138, B1 => l076_n_211, B2 => l076_n_126, C => l076_n_236, Z => l076_n_240);
  l076_g12418 : OAI32D0BWP7T port map(A1 => l076_n_26, A2 => l076_n_61, A3 => l076_n_221, B1 => l076_n_95, B2 => l076_n_223, ZN => b10);
  l076_g12419 : AOI211XD0BWP7T port map(A1 => l076_n_198, A2 => l076_n_70, B => l076_n_231, C => l076_n_225, ZN => l076_n_238);
  l076_g12420 : ND3D0BWP7T port map(A1 => l076_n_219, A2 => l076_n_210, A3 => l076_n_197, ZN => enable10);
  l076_g12421 : OAI211D1BWP7T port map(A1 => l076_n_84, A2 => l076_n_203, B => l076_n_218, C => l076_n_226, ZN => l076_n_236);
  l076_g12422 : ND4D0BWP7T port map(A1 => l076_n_215, A2 => l076_n_186, A3 => l076_n_180, A4 => l076_n_164, ZN => l076_n_235);
  l076_g12423 : OAI211D1BWP7T port map(A1 => l076_n_171, A2 => l076_n_223, B => l076_n_220, C => l076_n_206, ZN => l076_n_234);
  l076_g12424 : AOI22D0BWP7T port map(A1 => l076_n_211, A2 => l076_n_156, B1 => l076_n_216, B2 => l076_n_160, ZN => l076_n_233);
  l076_g12425 : AOI31D0BWP7T port map(A1 => l076_n_129, A2 => l076_n_131, A3 => l076_n_61, B => l076_n_229, ZN => l076_n_232);
  l076_g12426 : AOI21D0BWP7T port map(A1 => l076_n_131, A2 => l076_n_71, B => l076_n_224, ZN => l076_n_231);
  l076_g12427 : OAI21D0BWP7T port map(A1 => l076_n_132, A2 => l076_n_91, B => l076_n_222, ZN => l076_n_230);
  l076_g12428 : AOI21D0BWP7T port map(A1 => l076_n_209, A2 => l076_n_149, B => l076_n_195, ZN => l076_n_229);
  l076_g12429 : IAO21D0BWP7T port map(A1 => l076_n_152, A2 => l076_n_70, B => l076_n_212, ZN => l076_n_228);
  l076_g12430 : OAI31D0BWP7T port map(A1 => l076_n_75, A2 => l076_n_91, A3 => l076_n_111, B => l076_n_213, ZN => l076_n_227);
  l076_g12431 : OAI21D0BWP7T port map(A1 => l076_n_132, A2 => l076_n_138, B => l076_n_213, ZN => l076_n_226);
  l076_g12432 : AOI21D0BWP7T port map(A1 => l076_n_101, A2 => l076_n_69, B => l076_n_212, ZN => l076_n_225);
  l076_g12433 : CKND1BWP7T port map(I => l076_n_222, ZN => l076_n_223);
  l076_g12434 : OAI21D0BWP7T port map(A1 => l076_n_90, A2 => l076_n_55, B => l076_n_217, ZN => l076_n_220);
  l076_g12435 : AOI22D0BWP7T port map(A1 => l076_n_204, A2 => l076_n_192, B1 => l076_n_202, B2 => l076_n_177, ZN => l076_n_219);
  l076_g12436 : OAI21D0BWP7T port map(A1 => l076_n_92, A2 => l076_n_64, B => l076_n_216, ZN => l076_n_218);
  l076_g12437 : AOI22D0BWP7T port map(A1 => l076_n_208, A2 => l076_n_150, B1 => l076_n_209, B2 => l076_n_4, ZN => l076_n_224);
  l076_g12438 : OAI32D1BWP7T port map(A1 => l076_n_117, A2 => l076_n_134, A3 => l076_n_197, B1 => l076_n_157, B2 => l076_n_207, ZN => l076_n_222);
  l076_g12439 : AOI22D0BWP7T port map(A1 => l076_n_209, A2 => l076_n_6, B1 => l076_n_208, B2 => l076_n_151, ZN => l076_n_221);
  l076_g12440 : AOI211D1BWP7T port map(A1 => l076_n_127, A2 => l076_n_56, B => l076_n_196, C => l076_n_187, ZN => l076_n_215);
  l076_g12441 : OAI22D0BWP7T port map(A1 => l076_n_199, A2 => l076_n_170, B1 => l076_n_193, B2 => l076_n_180, ZN => l076_n_217);
  l076_g12442 : IOA21D1BWP7T port map(A1 => l076_n_202, A2 => l076_n_166, B => l076_n_210, ZN => l076_n_216);
  l076_g12443 : MOAI22D0BWP7T port map(A1 => l076_n_199, A2 => l076_n_164, B1 => l076_n_202, B2 => l076_n_165, ZN => l076_n_214);
  l076_g12444 : MOAI22D0BWP7T port map(A1 => l076_n_199, A2 => l076_n_167, B1 => l076_n_202, B2 => l076_n_168, ZN => l076_n_213);
  l076_g12445 : MAOI22D0BWP7T port map(A1 => l076_n_200, A2 => l076_n_165, B1 => l076_n_201, B2 => l076_n_164, ZN => l076_n_212);
  l076_g12446 : MOAI22D0BWP7T port map(A1 => l076_n_193, A2 => l076_n_186, B1 => l076_n_200, B2 => l076_n_166, ZN => l076_n_211);
  l076_g12447 : INVD0BWP7T port map(I => l076_n_208, ZN => l076_n_207);
  l076_g12448 : ND2D1BWP7T port map(A1 => l076_n_200, A2 => l076_n_148, ZN => l076_n_210);
  l076_g12449 : NR2D1BWP7T port map(A1 => l076_n_197, A2 => l076_n_112, ZN => l076_n_209);
  l076_g12450 : NR2D1BWP7T port map(A1 => l076_n_197, A2 => l076_n_113, ZN => l076_n_208);
  l076_g12451 : OAI21D0BWP7T port map(A1 => l076_n_130, A2 => l076_n_75, B => l076_n_198, ZN => l076_n_206);
  l076_g12452 : AOI21D0BWP7T port map(A1 => l076_n_142, A2 => l076_n_80, B => l076_n_203, ZN => l076_n_205);
  l076_g12453 : ND4D0BWP7T port map(A1 => l076_n_194, A2 => l076_n_189, A3 => l076_n_3, A4 => l076_n_181, ZN => l076_n_204);
  l076_g12454 : INVD0BWP7T port map(I => l076_n_202, ZN => l076_n_201);
  l076_g12455 : INVD0BWP7T port map(I => l076_n_200, ZN => l076_n_199);
  l076_g12456 : CKND2D1BWP7T port map(A1 => l076_n_192, A2 => l076_n_187, ZN => l076_n_203);
  l076_g12457 : NR2D1BWP7T port map(A1 => l076_n_193, A2 => l076_n_184, ZN => l076_n_202);
  l076_g12458 : NR2D1BWP7T port map(A1 => l076_n_193, A2 => l076_n_5, ZN => l076_n_200);
  l076_g12459 : OA31D1BWP7T port map(A1 => l076_n_119, A2 => l076_n_147, A3 => l076_n_174, B => l076_n_194, Z => l076_n_196);
  l076_g12460 : NR4D0BWP7T port map(A1 => l076_n_193, A2 => l076_n_172, A3 => l076_n_163, A4 => l076_n_43, ZN => l076_n_195);
  l076_g12461 : AOI21D0BWP7T port map(A1 => l076_n_3, A2 => l076_n_181, B => l076_n_193, ZN => l076_n_198);
  l076_g12462 : ND3D0BWP7T port map(A1 => l076_n_192, A2 => l076_n_175, A3 => l076_n_120, ZN => l076_n_197);
  l076_g12463 : INR2XD0BWP7T port map(A1 => l076_n_186, B1 => l076_n_191, ZN => l076_n_194);
  l076_g12464 : INVD1BWP7T port map(I => l076_n_193, ZN => l076_n_192);
  l076_g12465 : OAI221D0BWP7T port map(A1 => l076_n_173, A2 => l076_n_141, B1 => l076_n_30, B2 => l076_n_21, C => l076_n_190, ZN => l076_n_193);
  l076_g12466 : OAI221D0BWP7T port map(A1 => l076_n_5, A2 => l076_n_178, B1 => l076_n_170, B2 => l076_n_184, C => l076_n_180, ZN => l076_n_191);
  l076_g12467 : AOI221D0BWP7T port map(A1 => l076_n_9, A2 => x_enemy6(8), B1 => l076_n_51, B2 => l076_n_18, C => l076_n_185, ZN => l076_n_190);
  l076_g12468 : IAO21D0BWP7T port map(A1 => l076_n_184, A2 => l076_n_182, B => l076_n_188, ZN => l076_n_189);
  l076_g12469 : AOI21D0BWP7T port map(A1 => l076_n_182, A2 => l076_n_170, B => l076_n_5, ZN => l076_n_188);
  l076_g12470 : OAI22D0BWP7T port map(A1 => l076_n_184, A2 => l076_n_167, B1 => l076_n_5, B2 => l076_n_169, ZN => l076_n_187);
  l076_g12471 : IND2D1BWP7T port map(A1 => l076_n_184, B1 => l076_n_148, ZN => l076_n_186);
  l076_g12472 : AO21D0BWP7T port map(A1 => l076_n_21, A2 => l076_n_30, B => l076_n_179, Z => l076_n_185);
  l076_g12474 : NR3D0BWP7T port map(A1 => l076_n_162, A2 => l076_n_90, A3 => l076_n_64, ZN => l076_n_183);
  l076_g12476 : ND2D1BWP7T port map(A1 => l076_n_176, A2 => l076_n_118, ZN => l076_n_184);
  l076_g12477 : MOAI22D0BWP7T port map(A1 => l076_n_51, A2 => l076_n_18, B1 => l076_n_159, B2 => l076_n_141, ZN => l076_n_179);
  l076_g12478 : INR3D0BWP7T port map(A1 => l076_n_167, B1 => l076_n_165, B2 => l076_n_166, ZN => l076_n_182);
  l076_g12479 : ND4D0BWP7T port map(A1 => l076_n_1, A2 => l076_n_154, A3 => l076_n_145, A4 => l076_n_43, ZN => l076_n_181);
  l076_g12480 : IND3D1BWP7T port map(A1 => l076_n_147, B1 => l076_n_119, B2 => l076_n_176, ZN => l076_n_180);
  l076_g12481 : CKND1BWP7T port map(I => l076_n_177, ZN => l076_n_178);
  l076_g12482 : INVD0BWP7T port map(I => l076_n_175, ZN => l076_n_174);
  l076_g12483 : ND2D1BWP7T port map(A1 => l076_n_169, A2 => l076_n_164, ZN => l076_n_177);
  l076_g12484 : AOI211XD0BWP7T port map(A1 => l076_n_46, A2 => l076_n_31, B => l076_n_163, C => l076_n_100, ZN => l076_n_176);
  l076_g12485 : AOI211XD0BWP7T port map(A1 => l076_n_46, A2 => l076_n_25, B => l076_n_163, C => l076_n_99, ZN => l076_n_175);
  l076_g12486 : AOI221D0BWP7T port map(A1 => l076_n_106, A2 => l076_n_16, B1 => l076_n_49, B2 => l076_n_103, C => l076_n_158, ZN => l076_n_173);
  l076_g12487 : AOI22D0BWP7T port map(A1 => l076_n_1, A2 => y(4), B1 => l076_n_153, B2 => l076_n_41, ZN => l076_n_172);
  l076_g12488 : INR4D0BWP7T port map(A1 => l076_n_95, B1 => l076_n_93, B2 => l076_n_132, B3 => l076_n_146, ZN => l076_n_171);
  l076_g12489 : INVD0BWP7T port map(I => l076_n_169, ZN => l076_n_168);
  l076_g12490 : ND2D1BWP7T port map(A1 => l076_n_149, A2 => l076_n_112, ZN => l076_n_170);
  l076_g12491 : ND2D1BWP7T port map(A1 => l076_n_4, A2 => l076_n_112, ZN => l076_n_169);
  l076_g12492 : ND2D1BWP7T port map(A1 => l076_n_150, A2 => l076_n_113, ZN => l076_n_167);
  l076_g12493 : INR2D1BWP7T port map(A1 => l076_n_113, B1 => l076_n_157, ZN => l076_n_166);
  l076_g12494 : AN2D1BWP7T port map(A1 => l076_n_6, A2 => l076_n_112, Z => l076_n_165);
  l076_g12495 : ND2D1BWP7T port map(A1 => l076_n_151, A2 => l076_n_113, ZN => l076_n_164);
  l076_g12496 : IND4D0BWP7T port map(A1 => l076_n_70, B1 => l076_n_71, B2 => l076_n_101, B3 => l076_n_115, ZN => l076_n_162);
  l076_g12497 : ND4D0BWP7T port map(A1 => l076_n_128, A2 => l076_n_94, A3 => l076_n_69, A4 => l076_n_60, ZN => l076_n_161);
  l076_g12498 : IND4D0BWP7T port map(A1 => l076_n_75, B1 => l076_n_69, B2 => l076_n_76, B3 => l076_n_123, ZN => l076_n_160);
  l076_g12499 : OAI222D0BWP7T port map(A1 => l076_n_144, A2 => l076_n_137, B1 => l076_n_97, B2 => l076_n_136, C1 => l076_n_103, C2 => l076_n_104, ZN => l076_n_159);
  l076_g12500 : MOAI22D0BWP7T port map(A1 => l076_n_143, A2 => l076_n_135, B1 => l076_n_137, B2 => l076_n_105, ZN => l076_n_158);
  l076_g12501 : ND3D0BWP7T port map(A1 => l076_n_139, A2 => l076_n_145, A3 => l076_n_140, ZN => l076_n_163);
  l076_g12502 : OAI211D1BWP7T port map(A1 => l076_n_14, A2 => l076_n_56, B => l076_n_142, C => l076_n_88, ZN => l076_n_156);
  l076_g12503 : INR3D0BWP7T port map(A1 => l076_n_115, B1 => l076_n_92, B2 => l076_n_124, ZN => l076_n_155);
  l076_g12504 : AOI211D1BWP7T port map(A1 => l076_n_48, A2 => y(5), B => l076_n_122, C => l076_n_107, ZN => l076_n_154);
  l076_g12505 : NR3D0BWP7T port map(A1 => l076_n_133, A2 => l076_n_46, A3 => y(4), ZN => l076_n_153);
  l076_g12506 : AO211D0BWP7T port map(A1 => l076_n_59, A2 => l076_n_12, B => l076_n_146, C => l076_n_85, Z => l076_n_152);
  l076_g12507 : ND3D0BWP7T port map(A1 => l076_n_114, A2 => l076_n_109, A3 => l076_n_45, ZN => l076_n_157);
  l076_g12510 : NR3D0BWP7T port map(A1 => l076_n_116, A2 => l076_n_45, A3 => l076_n_47, ZN => l076_n_151);
  l076_g12512 : NR3D0BWP7T port map(A1 => l076_n_121, A2 => l076_n_114, A3 => l076_n_44, ZN => l076_n_150);
  l076_g12513 : AN4D1BWP7T port map(A1 => l076_n_114, A2 => l076_n_2, A3 => l076_n_108, A4 => l076_n_45, Z => l076_n_149);
  l076_g12514 : INR2D1BWP7T port map(A1 => l076_n_117, B1 => l076_n_134, ZN => l076_n_148);
  l076_g12515 : OR2D1BWP7T port map(A1 => l076_n_133, A2 => l076_n_41, Z => l076_n_147);
  l076_g12516 : ND2D1BWP7T port map(A1 => l076_n_131, A2 => l076_n_94, ZN => l076_n_146);
  l076_g12517 : AOI211XD0BWP7T port map(A1 => l076_n_53, A2 => l076_n_34, B => l076_n_89, C => l076_n_110, ZN => l076_n_145);
  l076_g12518 : CKND1BWP7T port map(I => l076_n_143, ZN => l076_n_144);
  l076_g12519 : AOI22D0BWP7T port map(A1 => l076_n_98, A2 => y(5), B1 => l076_n_82, B2 => y_enemy6(5), ZN => l076_n_140);
  l076_g12520 : NR2XD0BWP7T port map(A1 => l076_n_122, A2 => l076_n_107, ZN => l076_n_139);
  l076_g12521 : MAOI222D1BWP7T port map(A => l076_n_87, B => x(2), C => x_enemy6(2), ZN => l076_n_143);
  l076_g12522 : NR3D0BWP7T port map(A1 => l076_n_96, A2 => l076_n_90, A3 => l076_n_68, ZN => l076_n_142);
  l076_g12523 : OAI21D0BWP7T port map(A1 => l076_n_106, A2 => l076_n_15, B => l076_n_104, ZN => l076_n_141);
  l076_g12524 : CKND1BWP7T port map(I => l076_n_135, ZN => l076_n_136);
  l076_g12525 : INVD0BWP7T port map(I => l076_n_131, ZN => l076_n_130);
  l076_g12526 : AOI211XD0BWP7T port map(A1 => l076_n_59, A2 => l076_n_26, B => l076_n_96, C => l076_n_79, ZN => l076_n_129);
  l076_g12527 : OAI21D0BWP7T port map(A1 => l076_n_73, A2 => l076_n_58, B => draw_count10(1), ZN => l076_n_128);
  l076_g12528 : AOI221D0BWP7T port map(A1 => l076_n_58, A2 => l076_n_27, B1 => l076_n_62, B2 => draw_count10(0), C => l076_n_77, ZN => l076_n_127);
  l076_g12529 : AO221D0BWP7T port map(A1 => l076_n_65, A2 => l076_n_64, B1 => l076_n_66, B2 => l076_n_28, C => l076_n_93, Z => l076_n_126);
  l076_g12530 : OA211D0BWP7T port map(A1 => l076_n_26, A2 => l076_n_60, B => l076_n_101, C => l076_n_78, Z => l076_n_125);
  l076_g12531 : OAI211D1BWP7T port map(A1 => l076_n_12, A2 => l076_n_56, B => l076_n_80, C => l076_n_74, ZN => l076_n_124);
  l076_g12532 : AOI21D0BWP7T port map(A1 => l076_n_59, A2 => l076_n_27, B => l076_n_86, ZN => l076_n_123);
  l076_g12533 : AO21D0BWP7T port map(A1 => l076_n_66, A2 => l076_n_65, B => l076_n_93, Z => l076_n_138);
  l076_g12534 : OAI22D0BWP7T port map(A1 => l076_n_67, A2 => l076_n_17, B1 => l076_n_50, B2 => x(2), ZN => l076_n_137);
  l076_g12535 : IOA21D1BWP7T port map(A1 => l076_n_50, A2 => x(2), B => l076_n_105, ZN => l076_n_135);
  l076_g12536 : ND2D1BWP7T port map(A1 => l076_n_102, A2 => l076_n_42, ZN => l076_n_134);
  l076_g12537 : ND2D1BWP7T port map(A1 => l076_n_102, A2 => l076_n_83, ZN => l076_n_133);
  l076_g12538 : IND2D1BWP7T port map(A1 => l076_n_92, B1 => l076_n_69, ZN => l076_n_132);
  l076_g12539 : INR2XD0BWP7T port map(A1 => l076_n_60, B1 => l076_n_90, ZN => l076_n_131);
  l076_g12544 : OAI22D0BWP7T port map(A1 => l076_n_52, A2 => l076_n_29, B1 => l076_n_48, B2 => y(5), ZN => l076_n_122);
  l076_g12545 : MOAI22D0BWP7T port map(A1 => l076_n_60, A2 => draw_count10(1), B1 => l076_n_73, B2 => l076_n_65, ZN => l076_n_111);
  l076_g12546 : MOAI22D0BWP7T port map(A1 => l076_n_20, A2 => y(9), B1 => l076_n_20, B2 => y(9), ZN => l076_n_110);
  l076_g12547 : MAOI22D0BWP7T port map(A1 => l076_n_83, A2 => l076_n_35, B1 => l076_n_83, B2 => l076_n_35, ZN => l076_n_121);
  l076_g12548 : MAOI22D0BWP7T port map(A1 => l076_n_43, A2 => l076_n_36, B1 => l076_n_43, B2 => l076_n_36, ZN => l076_n_120);
  l076_g12549 : MAOI22D0BWP7T port map(A1 => l076_n_43, A2 => y(3), B1 => l076_n_43, B2 => y(3), ZN => l076_n_119);
  l076_g12550 : MAOI22D0BWP7T port map(A1 => l076_n_43, A2 => l076_n_19, B1 => l076_n_43, B2 => l076_n_19, ZN => l076_n_118);
  l076_g12551 : MAOI22D0BWP7T port map(A1 => l076_n_81, A2 => y(2), B1 => l076_n_81, B2 => y(2), ZN => l076_n_117);
  l076_g12552 : ND2D1BWP7T port map(A1 => l076_n_2, A2 => l076_n_108, ZN => l076_n_109);
  l076_g12553 : MAOI22D0BWP7T port map(A1 => l076_n_42, A2 => y(1), B1 => l076_n_42, B2 => y(1), ZN => l076_n_116);
  l076_g12554 : INR3D0BWP7T port map(A1 => l076_n_78, B1 => l076_n_62, B2 => l076_n_77, ZN => l076_n_115);
  l076_g12555 : MOAI22D0BWP7T port map(A1 => l076_n_47, A2 => y(0), B1 => l076_n_47, B2 => y(0), ZN => l076_n_114);
  l076_g12556 : MAOI22D0BWP7T port map(A1 => l076_n_41, A2 => l076_n_22, B1 => l076_n_41, B2 => l076_n_22, ZN => l076_n_113);
  l076_g12557 : MOAI22D0BWP7T port map(A1 => l076_n_41, A2 => l076_n_24, B1 => l076_n_41, B2 => l076_n_24, ZN => l076_n_112);
  l076_g12558 : NR2XD0BWP7T port map(A1 => l076_n_46, A2 => l076_n_31, ZN => l076_n_100);
  l076_g12559 : NR2D0BWP7T port map(A1 => l076_n_46, A2 => l076_n_25, ZN => l076_n_99);
  l076_g12560 : ND2D1BWP7T port map(A1 => l076_n_83, A2 => l076_n_32, ZN => l076_n_108);
  l076_g12561 : AN2D1BWP7T port map(A1 => l076_n_52, A2 => l076_n_29, Z => l076_n_107);
  l076_g12563 : NR2D0BWP7T port map(A1 => l076_n_82, A2 => y_enemy6(5), ZN => l076_n_98);
  l076_g12564 : CKAN2D1BWP7T port map(A1 => l076_n_49, A2 => l076_n_39, Z => l076_n_106);
  l076_g12565 : ND2D1BWP7T port map(A1 => l076_n_67, A2 => l076_n_17, ZN => l076_n_105);
  l076_g12566 : OR2D1BWP7T port map(A1 => l076_n_49, A2 => l076_n_16, Z => l076_n_104);
  l076_g12567 : NR2XD0BWP7T port map(A1 => l076_n_67, A2 => l076_n_17, ZN => l076_n_97);
  l076_g12568 : CKAN2D1BWP7T port map(A1 => l076_n_15, A2 => l076_n_39, Z => l076_n_103);
  l076_g12569 : INR2D1BWP7T port map(A1 => l076_n_47, B1 => l076_n_45, ZN => l076_n_102);
  l076_g12570 : NR2XD0BWP7T port map(A1 => l076_n_72, A2 => l076_n_79, ZN => l076_n_101);
  l076_g12571 : NR2D0BWP7T port map(A1 => l076_n_53, A2 => l076_n_34, ZN => l076_n_89);
  l076_g12572 : AOI22D0BWP7T port map(A1 => l076_n_59, A2 => l076_n_13, B1 => l076_n_62, B2 => l076_n_26, ZN => l076_n_88);
  l076_g12573 : AOI22D0BWP7T port map(A1 => l076_n_54, A2 => x(0), B1 => x(1), B2 => l076_n_10, ZN => l076_n_87);
  l076_g12574 : AOI21D0BWP7T port map(A1 => l076_n_57, A2 => l076_n_60, B => draw_count10(1), ZN => l076_n_86);
  l076_g12575 : OA21D0BWP7T port map(A1 => l076_n_58, A2 => l076_n_55, B => l076_n_26, Z => l076_n_85);
  l076_g12576 : AOI21D0BWP7T port map(A1 => l076_n_58, A2 => l076_n_26, B => l076_n_63, ZN => l076_n_84);
  l076_g12577 : OAI21D0BWP7T port map(A1 => l076_n_56, A2 => draw_count10(1), B => l076_n_74, ZN => l076_n_96);
  l076_g12578 : AOI21D0BWP7T port map(A1 => l076_n_62, A2 => l076_n_12, B => l076_n_59, ZN => l076_n_95);
  l076_g12579 : OAI21D0BWP7T port map(A1 => l076_n_63, A2 => l076_n_55, B => l076_n_13, ZN => l076_n_94);
  l076_g12580 : MOAI22D0BWP7T port map(A1 => l076_n_0, A2 => l076_n_27, B1 => l076_n_66, B2 => l076_n_13, ZN => l076_n_93);
  l076_g12581 : AO21D0BWP7T port map(A1 => l076_n_64, A2 => l076_n_27, B => l076_n_72, Z => l076_n_92);
  l076_g12582 : IOA21D1BWP7T port map(A1 => l076_n_58, A2 => l076_n_12, B => l076_n_76, ZN => l076_n_91);
  l076_g12583 : OAI22D0BWP7T port map(A1 => l076_n_57, A2 => l076_n_12, B1 => l076_n_60, B2 => l076_n_27, ZN => l076_n_90);
  l076_g12584 : INVD1BWP7T port map(I => l076_n_42, ZN => l076_n_83);
  l076_g12586 : INVD0BWP7T port map(I => l076_n_48, ZN => l076_n_82);
  l076_g12587 : INVD0BWP7T port map(I => l076_n_41, ZN => l076_n_81);
  l076_g12588 : ND2D1BWP7T port map(A1 => l076_n_59, A2 => draw_count10(1), ZN => l076_n_80);
  l076_g12589 : NR2D1BWP7T port map(A1 => l076_n_0, A2 => draw_count10(1), ZN => l076_n_79);
  l076_g12590 : IND2D0BWP7T port map(A1 => l076_n_14, B1 => l076_n_63, ZN => l076_n_78);
  l076_g12591 : INR2D1BWP7T port map(A1 => l076_n_59, B1 => draw_count10(1), ZN => l076_n_77);
  l076_g12592 : CKND2D0BWP7T port map(A1 => l076_n_63, A2 => l076_n_13, ZN => l076_n_76);
  l076_g12593 : NR2D0BWP7T port map(A1 => l076_n_56, A2 => l076_n_7, ZN => l076_n_75);
  l076_g12594 : NR2D0BWP7T port map(A1 => l076_n_60, A2 => l076_n_14, ZN => l076_n_68);
  l076_g12595 : CKND2D1BWP7T port map(A1 => l076_n_58, A2 => l076_n_65, ZN => l076_n_74);
  l076_g12596 : IND2D1BWP7T port map(A1 => l076_n_59, B1 => l076_n_61, ZN => l076_n_73);
  l076_g12597 : AN2D0BWP7T port map(A1 => l076_n_63, A2 => l076_n_26, Z => l076_n_72);
  l076_g12598 : ND2D1BWP7T port map(A1 => l076_n_55, A2 => l076_n_12, ZN => l076_n_71);
  l076_g12599 : INR2D1BWP7T port map(A1 => l076_n_28, B1 => l076_n_57, ZN => l076_n_70);
  l076_g12600 : ND2D1BWP7T port map(A1 => l076_n_63, A2 => l076_n_65, ZN => l076_n_69);
  l076_g12601 : INVD1BWP7T port map(I => l076_n_0, ZN => l076_n_64);
  l076_g12602 : INVD0BWP7T port map(I => l076_n_62, ZN => l076_n_61);
  l076_g12603 : INVD0BWP7T port map(I => l076_n_58, ZN => l076_n_57);
  l076_g12604 : INVD1BWP7T port map(I => l076_n_56, ZN => l076_n_55);
  l076_g12605 : IAO21D0BWP7T port map(A1 => x(1), A2 => l076_n_10, B => x_enemy6(0), ZN => l076_n_54);
  l076_g12606 : AO21D0BWP7T port map(A1 => x(4), A2 => l076_n_11, B => l076_n_15, Z => l076_n_67);
  l076_g12607 : INR2D1BWP7T port map(A1 => draw_count10(3), B1 => l076_n_33, ZN => l076_n_66);
  l076_g12608 : IND2D1BWP7T port map(A1 => l076_n_28, B1 => l076_n_14, ZN => l076_n_65);
  l076_g12610 : NR2D1BWP7T port map(A1 => l076_n_33, A2 => draw_count10(3), ZN => l076_n_63);
  l076_g12611 : INR2D1BWP7T port map(A1 => l076_n_23, B1 => draw_count10(3), ZN => l076_n_62);
  l076_g12612 : ND2D1BWP7T port map(A1 => l076_n_37, A2 => draw_count10(3), ZN => l076_n_60);
  l076_g12613 : NR2D1BWP7T port map(A1 => l076_n_38, A2 => draw_count10(3), ZN => l076_n_59);
  l076_g12614 : NR2D1BWP7T port map(A1 => l076_n_40, A2 => draw_count10(3), ZN => l076_n_58);
  l076_g12615 : ND2D1BWP7T port map(A1 => l076_n_23, A2 => draw_count10(3), ZN => l076_n_56);
  l076_g12617 : INVD0BWP7T port map(I => l076_n_45, ZN => l076_n_44);
  l076_g12618 : MOAI22D0BWP7T port map(A1 => y(8), A2 => y_enemy6(8), B1 => y(8), B2 => y_enemy6(8), ZN => l076_n_53);
  l076_g12619 : MAOI22D0BWP7T port map(A1 => y(7), A2 => y_enemy6(7), B1 => y(7), B2 => y_enemy6(7), ZN => l076_n_52);
  l076_g12620 : MOAI22D0BWP7T port map(A1 => x(7), A2 => x_enemy6(7), B1 => x(7), B2 => x_enemy6(7), ZN => l076_n_51);
  l076_g12621 : MAOI22D0BWP7T port map(A1 => x(3), A2 => x_enemy6(3), B1 => x(3), B2 => x_enemy6(3), ZN => l076_n_50);
  l076_g12622 : MAOI22D0BWP7T port map(A1 => x(6), A2 => x_enemy6(6), B1 => x(6), B2 => x_enemy6(6), ZN => l076_n_49);
  l076_g12623 : OAI21D0BWP7T port map(A1 => l076_n_8, A2 => y_enemy6(6), B => l076_n_29, ZN => l076_n_48);
  l076_g12624 : MOAI22D0BWP7T port map(A1 => y(1), A2 => y_enemy6(1), B1 => y(1), B2 => y_enemy6(1), ZN => l076_n_47);
  l076_g12625 : MAOI22D0BWP7T port map(A1 => y(5), A2 => y_enemy6(5), B1 => y(5), B2 => y_enemy6(5), ZN => l076_n_46);
  l076_g12626 : MAOI22D0BWP7T port map(A1 => y(0), A2 => y_enemy6(0), B1 => y(0), B2 => y_enemy6(0), ZN => l076_n_45);
  l076_g12627 : MOAI22D0BWP7T port map(A1 => y(4), A2 => y_enemy6(4), B1 => y(4), B2 => y_enemy6(4), ZN => l076_n_43);
  l076_g12628 : MAOI22D0BWP7T port map(A1 => y(2), A2 => y_enemy6(2), B1 => y(2), B2 => y_enemy6(2), ZN => l076_n_42);
  l076_g12629 : MOAI22D0BWP7T port map(A1 => y(3), A2 => y_enemy6(3), B1 => y(3), B2 => y_enemy6(3), ZN => l076_n_41);
  l076_g12631 : CKND1BWP7T port map(I => l076_n_37, ZN => l076_n_38);
  l076_g12632 : INVD1BWP7T port map(I => l076_n_27, ZN => l076_n_26);
  l076_g12633 : IND2D1BWP7T port map(A1 => draw_count10(2), B1 => draw_count10(4), ZN => l076_n_40);
  l076_g12634 : IND2D1BWP7T port map(A1 => x_enemy6(5), B1 => x(5), ZN => l076_n_39);
  l076_g12635 : INR2D1BWP7T port map(A1 => draw_count10(2), B1 => draw_count10(4), ZN => l076_n_37);
  l076_g12636 : IND2D0BWP7T port map(A1 => y_enemy6(3), B1 => y(3), ZN => l076_n_36);
  l076_g12637 : IND2D0BWP7T port map(A1 => y_enemy6(1), B1 => y(1), ZN => l076_n_35);
  l076_g12638 : INR2XD0BWP7T port map(A1 => y_enemy6(7), B1 => y(7), ZN => l076_n_34);
  l076_g12639 : ND2D1BWP7T port map(A1 => draw_count10(2), A2 => draw_count10(4), ZN => l076_n_33);
  l076_g12640 : INR2XD0BWP7T port map(A1 => y_enemy6(1), B1 => y(1), ZN => l076_n_32);
  l076_g12641 : IND2D1BWP7T port map(A1 => y_enemy6(4), B1 => y(4), ZN => l076_n_31);
  l076_g12642 : IND2D1BWP7T port map(A1 => x(7), B1 => x_enemy6(7), ZN => l076_n_30);
  l076_g12643 : ND2D1BWP7T port map(A1 => l076_n_8, A2 => y_enemy6(6), ZN => l076_n_29);
  l076_g12644 : INR2D1BWP7T port map(A1 => draw_count10(0), B1 => draw_count10(1), ZN => l076_n_28);
  l076_g12645 : CKND2D1BWP7T port map(A1 => draw_count10(1), A2 => draw_count10(0), ZN => l076_n_27);
  l076_g12646 : INVD1BWP7T port map(I => l076_n_13, ZN => l076_n_12);
  l076_g12647 : INR2XD0BWP7T port map(A1 => y_enemy6(4), B1 => y(4), ZN => l076_n_25);
  l076_g12648 : IND2D1BWP7T port map(A1 => y(2), B1 => y_enemy6(2), ZN => l076_n_24);
  l076_g12649 : NR2D0BWP7T port map(A1 => draw_count10(2), A2 => draw_count10(4), ZN => l076_n_23);
  l076_g12650 : IND2D1BWP7T port map(A1 => y_enemy6(2), B1 => y(2), ZN => l076_n_22);
  l076_g12651 : NR2D0BWP7T port map(A1 => l076_n_9, A2 => x_enemy6(8), ZN => l076_n_21);
  l076_g12652 : IND2D1BWP7T port map(A1 => y(8), B1 => y_enemy6(8), ZN => l076_n_20);
  l076_g12653 : IND2D1BWP7T port map(A1 => y(3), B1 => y_enemy6(3), ZN => l076_n_19);
  l076_g12654 : IND2D1BWP7T port map(A1 => x_enemy6(6), B1 => x(6), ZN => l076_n_18);
  l076_g12655 : IND2D1BWP7T port map(A1 => x(3), B1 => x_enemy6(3), ZN => l076_n_17);
  l076_g12656 : INR2XD0BWP7T port map(A1 => x_enemy6(5), B1 => x(5), ZN => l076_n_16);
  l076_g12657 : NR2D0BWP7T port map(A1 => x(4), A2 => l076_n_11, ZN => l076_n_15);
  l076_g12658 : IND2D1BWP7T port map(A1 => draw_count10(0), B1 => draw_count10(1), ZN => l076_n_14);
  l076_g12659 : NR2D0BWP7T port map(A1 => draw_count10(1), A2 => draw_count10(0), ZN => l076_n_13);
  l076_g12660 : CKND1BWP7T port map(I => x_enemy6(4), ZN => l076_n_11);
  l076_g12661 : INVD0BWP7T port map(I => x_enemy6(1), ZN => l076_n_10);
  l076_g12662 : CKND1BWP7T port map(I => x(8), ZN => l076_n_9);
  l076_g12663 : CKND1BWP7T port map(I => y(6), ZN => l076_n_8);
  l076_g12664 : INVD0BWP7T port map(I => draw_count10(1), ZN => l076_n_7);
  l076_g2 : INR3D0BWP7T port map(A1 => l076_n_121, B1 => l076_n_114, B2 => l076_n_44, ZN => l076_n_6);
  l076_g12665 : IND2D1BWP7T port map(A1 => l076_n_118, B1 => l076_n_175, ZN => l076_n_5);
  l076_g12666 : INR3D0BWP7T port map(A1 => l076_n_116, B1 => l076_n_45, B2 => l076_n_47, ZN => l076_n_4);
  l076_g12667 : IIND4D0BWP7T port map(A1 => l076_n_120, A2 => l076_n_112, B1 => l076_n_149, B2 => l076_n_176, ZN => l076_n_3);
  l076_g12668 : IND2D1BWP7T port map(A1 => l076_n_32, B1 => l076_n_42, ZN => l076_n_2);
  l076_g12669 : INR3D0BWP7T port map(A1 => l076_n_46, B1 => l076_n_133, B2 => l076_n_81, ZN => l076_n_1);
  l076_g12670 : IND2D1BWP7T port map(A1 => l076_n_40, B1 => draw_count10(3), ZN => l076_n_0);
  l041_count_reg_2 : DFCNQD1BWP7T port map(CDN => l041_n_0, CP => clk, D => l041_n_6, Q => draw_count1(2));
  l041_g59 : CKAN2D1BWP7T port map(A1 => enable1, A2 => l041_n_5, Z => l041_n_6);
  l041_count_reg_1 : DFCNQD1BWP7T port map(CDN => l041_n_0, CP => clk, D => l041_n_4, Q => draw_count1(1));
  l041_g61 : MOAI22D0BWP7T port map(A1 => l041_n_1, A2 => draw_count1(2), B1 => l041_n_1, B2 => draw_count1(2), ZN => l041_n_5);
  l041_g62 : CKAN2D1BWP7T port map(A1 => enable1, A2 => l041_n_3, Z => l041_n_4);
  l041_count_reg_0 : DFCNQD1BWP7T port map(CDN => l041_n_0, CP => clk, D => l041_n_2, Q => draw_count1(0));
  l041_g64 : CKXOR2D1BWP7T port map(A1 => draw_count1(0), A2 => draw_count1(1), Z => l041_n_3);
  l041_g65 : INR2XD0BWP7T port map(A1 => enable1, B1 => draw_count1(0), ZN => l041_n_2);
  l041_g66 : ND2D1BWP7T port map(A1 => draw_count1(1), A2 => draw_count1(0), ZN => l041_n_1);
  l041_g67 : INVD0BWP7T port map(I => reset, ZN => l041_n_0);

end synthesised;
