configuration top_level_routed_cfg of top_level is
   for routed
   end for;
end top_level_routed_cfg;
