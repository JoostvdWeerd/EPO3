configuration bullet_behaviour_cfg of bullet is
   for behaviour
   end for;
end bullet_behaviour_cfg;
