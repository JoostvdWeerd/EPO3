configuration sync_behaviour_cfg of sync is
   for behaviour
   end for;
end sync_behaviour_cfg;
