library IEEE;
use IEEE.std_logic_1164.ALL;

entity display_tb is
end display_tb;

