configuration x_counter_behaviour_cfg of x_counter is
   for behaviour
   end for;
end x_counter_behaviour_cfg;
