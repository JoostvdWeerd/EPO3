configuration collision_behaviour_collision_cfg of collision is
   for behaviour_collision
   end for;
end collision_behaviour_collision_cfg;
