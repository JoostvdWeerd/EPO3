configuration display_routed_cfg of display is
   for routed
   end for;
end display_routed_cfg;
