configuration y_counter_behaviour_cfg of y_counter is
   for behaviour
   end for;
end y_counter_behaviour_cfg;
