configuration top_level_synthesised_cfg of top_level is
   for synthesised
   end for;
end top_level_synthesised_cfg;
