configuration counter_one_behaviour_counter_one_cfg of counter_one is
   for behaviour_counter_one
   end for;
end counter_one_behaviour_counter_one_cfg;
