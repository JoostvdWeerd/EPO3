configuration display_tb_behaviour_rou_cfg of display_tb is
   for behaviour
      for all: display use configuration work.display_routed_cfg;
      end for;
   end for;
end display_tb_behaviour_rou_cfg;
