configuration counter_two_behaviour_counter_two_cfg of counter_two is
   for behaviour_counter_two
   end for;
end counter_two_behaviour_counter_two_cfg;
